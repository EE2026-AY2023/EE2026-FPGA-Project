`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.03.2023 18:48:27
// Design Name: 
// Module Name: end_screen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

//explosion credits:https://www.reddit.com/r/PixelArt/comments/wvtxti/explosion_effect_from_a_series_of_vfx_im_working/
//<a href="https://www.freepik.com/free-vector/pixelated-trophy-card-with-lettering_29171430.htm">Image by gstudioimagen1</a> on Freepik
module ftb_end_loss_screen(
    input clock,
    input [6:0] x, y,
    output reg [15:0] oled_data = 0
    );
    always @(posedge clock) begin
        if ((y == 50 && x == 41)) oled_data <= 16'hfbef;
        else if ((y == 40 && x == 36)) oled_data <= 16'h58cd;
        else if ((y == 48 && x == 28) || (y == 50 && x == 30) || (y == 48 && x == 31) || (y == 50 && x == 33) || (y == 50 && x == 59) || (y == 49 && x == 61) || (y == 48 && x == 69)) oled_data <= 16'ha1ce;
        else if ((y == 19 && x == 58)) oled_data <= 16'h6817;
        else if ((y == 22 && x == 42) || (y == 22 && x == 52) || (y == 30 && x == 62)) oled_data <= 16'h29a9;
        else if ((y == 31 && x == 41)) oled_data <= 16'h1d99;
        else if ((y == 23 && x == 47)) oled_data <= 16'h12d5;
        else if ((y == 33 && x == 25) || (y == 41 && x == 73)) oled_data <= 16'h31a7;
        else if ((y == 46 && x == 62)) oled_data <= 16'hb517;
        else if ((y == 52 && x == 42)) oled_data <= 16'h79ed;
        else if ((y == 45 && x == 44)) oled_data <= 16'hac09;
        else if ((y == 51 && x == 44)) oled_data <= 16'hff7f;
        else if ((y == 30 && x == 45) || (y == 36 && x == 57)) oled_data <= 16'ha00a;
        else if ((y == 52 && x == 52)) oled_data <= 16'hc212;
        else if ((y == 36 && x == 31)) oled_data <= 16'h31cc;
        else if ((y == 44 && x == 43)) oled_data <= 16'hfbc0;
        else if ((y == 27 && x == 52)) oled_data <= 16'hf081;
        else if ((y == 32 && x == 37)) oled_data <= 16'h16be;
        else if ((y == 31 && x == 58)) oled_data <= 16'h490d;
        else if ((y == 31 && x == 71)) oled_data <= 16'h4838;
        else if ((y == 20 && x == 38) || (y == 19 && x == 41) || (y == 18 && x == 44) || (y == 18 && x == 45) || (y == 18 && x == 46) || (y == 18 && x == 52) || (y == 18 && x == 53) || (y == 19 && x == 56) || (y == 19 && x == 57) || (y == 20 && x == 60) || (y == 21 && x == 61)) oled_data <= 16'h6015;
        else if ((y == 35 && x == 40)) oled_data <= 16'hc2f1;
        else if ((y == 42 && x == 41) || (y == 38 && x == 49)) oled_data <= 16'hfc60;
        else if ((y == 37 && x == 39)) oled_data <= 16'hf980;
        else if ((y == 47 && x == 58)) oled_data <= 16'h16ff;
        else if ((y == 51 && x == 41)) oled_data <= 16'hd254;
        else if ((y == 47 && x == 24) || (y == 48 && x == 24) || (y == 47 && x == 25) || (y == 48 && x == 25) || (y == 45 && x == 26) || (y == 48 && x == 26) || (y == 49 && x == 26) || (y == 47 && x == 28) || (y == 50 && x == 28) || (y == 45 && x == 29) || (y == 48 && x == 29) || (y == 48 && x == 30) || (y == 49 && x == 30) || (y == 49 && x == 31) || (y == 50 && x == 31) || (y == 48 && x == 32) || (y == 50 && x == 32) || (y == 52 && x == 33) || (y == 52 && x == 34) || (y == 53 && x == 34) || (y == 49 && x == 35) || (y == 50 && x == 35) || (y == 51 && x == 35) || (y == 52 && x == 35) || (y == 53 && x == 35) || (y == 51 && x == 36) || (y == 52 && x == 36) || (y == 53 && x == 36) || (y == 52 && x == 37) || (y == 52 && x == 38) || (y == 52 && x == 39) || (y == 55 && x == 39) || (y == 53 && x == 40) || (y == 55 && x == 40) || (y == 53 && x == 41) || (y == 53 && x == 42) || (y == 54 && x == 44) || (y == 55 && x == 44) || (y == 54 && x == 45) || (y == 55 && x == 45) || (y == 54 && x == 46) || (y == 54 && x == 47) || (y == 56 && x == 47) || (y == 56 && x == 48) || (y == 56 && x == 49) || (y == 53 && x == 50) || (y == 54 && x == 50) || (y == 56 && x == 50) || (y == 54 && x == 51) || (y == 56 && x == 51) || (y == 54 && x == 52) || (y == 54 && x == 53) || (y == 55 && x == 53) || (y == 53 && x == 54) || (y == 53 && x == 55) || (y == 52 && x == 56) || (y == 53 && x == 56) || (y == 55 && x == 56) || (y == 52 && x == 57) || (y == 53 && x == 57) || (y == 54 && x == 57) || (y == 55 && x == 57) || (y == 52 && x == 58) || (y == 53 && x == 58) || (y == 54 && x == 58) || (y == 55 && x == 58) || (y == 51 && x == 59) || (y == 52 && x == 59) || (y == 53 && x == 59) || (y == 55 && x == 59) || (y == 50 && x == 60) || (y == 53 && x == 60) || (y == 55 && x == 60) || (y == 50 && x == 61) || (y == 52 && x == 61) || (y == 53 && x == 61) || (y == 52 && x == 62) || (y == 54 && x == 62) || (y == 52 && x == 63) || (y == 48 && x == 64) || (y == 51 && x == 64) || (y == 52 && x == 64) || (y == 44 && x == 65) || (y == 45 && x == 65) || (y == 47 && x == 65) || (y == 48 && x == 65) || (y == 49 && x == 65) || (y == 50 && x == 65) || (y == 51 && x == 65) || (y == 44 && x == 66) || (y == 45 && x == 66) || (y == 46 && x == 66) || (y == 47 && x == 66) || (y == 48 && x == 66) || (y == 50 && x == 66) || (y == 51 && x == 66) || (y == 52 && x == 66) || (y == 47 && x == 67) || (y == 49 && x == 67) || (y == 50 && x == 67) || (y == 51 && x == 67) || (y == 52 && x == 67) || (y == 46 && x == 68) || (y == 49 && x == 68) || (y == 51 && x == 68) || (y == 49 && x == 69) || (y == 43 && x == 70) || (y == 48 && x == 70) || (y == 42 && x == 71) || (y == 47 && x == 71) || (y == 41 && x == 72)) oled_data <= 16'h520b;
        else if ((y == 35 && x == 25) || (y == 36 && x == 25) || (y == 37 && x == 25) || (y == 44 && x == 25) || (y == 35 && x == 72) || (y == 43 && x == 72)) oled_data <= 16'h201f;
        else if ((y == 31 && x == 55)) oled_data <= 16'h8ad2;
        else if ((y == 38 && x == 29)) oled_data <= 16'h4992;
        else if ((y == 51 && x == 34)) oled_data <= 16'h91ce;
        else if ((y == 36 && x == 44) || (y == 43 && x == 54) || (y == 47 && x == 55)) oled_data <= 16'hfac0;
        else if ((y == 47 && x == 39) || (y == 48 && x == 39) || (y == 46 && x == 40) || (y == 47 && x == 40) || (y == 48 && x == 40) || (y == 49 && x == 40) || (y == 46 && x == 41) || (y == 49 && x == 41) || (y == 41 && x == 42) || (y == 48 && x == 42) || (y == 49 && x == 42) || (y == 40 && x == 43) || (y == 40 && x == 44) || (y == 43 && x == 44) || (y == 44 && x == 44) || (y == 38 && x == 45) || (y == 40 && x == 45) || (y == 42 && x == 45) || (y == 43 && x == 45) || (y == 44 && x == 45) || (y == 38 && x == 46) || (y == 39 && x == 46) || (y == 40 && x == 46) || (y == 42 && x == 46) || (y == 43 && x == 46) || (y == 44 && x == 46) || (y == 38 && x == 47) || (y == 39 && x == 47) || (y == 40 && x == 47) || (y == 42 && x == 47) || (y == 43 && x == 47) || (y == 39 && x == 48) || (y == 40 && x == 48) || (y == 42 && x == 48) || (y == 32 && x == 49) || (y == 40 && x == 49) || (y == 33 && x == 50) || (y == 38 && x == 50) || (y == 39 && x == 51) || (y == 43 && x == 51) || (y == 42 && x == 52) || (y == 43 && x == 52) || (y == 44 && x == 52) || (y == 42 && x == 53) || (y == 43 && x == 53) || (y == 44 && x == 53) || (y == 46 && x == 53) || (y == 47 && x == 53) || (y == 49 && x == 53) || (y == 47 && x == 54) || (y == 48 && x == 54) || (y == 49 && x == 54) || (y == 50 && x == 54) || (y == 49 && x == 55) || (y == 50 && x == 55)) oled_data <= 16'hfe60;
        else if ((y == 46 && x == 31)) oled_data <= 16'hd275;
        else if ((y == 31 && x == 26) || (y == 29 && x == 27) || (y == 19 && x == 42) || (y == 18 && x == 55) || (y == 19 && x == 55) || (y == 29 && x == 69)) oled_data <= 16'h29c7;
        else if ((y == 46 && x == 34)) oled_data <= 16'he276;
        else if ((y == 44 && x == 42)) oled_data <= 16'hfdc0;
        else if ((y == 32 && x == 38)) oled_data <= 16'hf7bf;
        else if ((y == 48 && x == 27) || (y == 49 && x == 27) || (y == 46 && x == 28) || (y == 49 && x == 28) || (y == 46 && x == 29) || (y == 49 && x == 29) || (y == 50 && x == 29) || (y == 44 && x == 32) || (y == 45 && x == 32) || (y == 46 && x == 32) || (y == 48 && x == 34) || (y == 47 && x == 36) || (y == 49 && x == 36) || (y == 50 && x == 36) || (y == 49 && x == 37) || (y == 50 && x == 37) || (y == 50 && x == 38) || (y == 51 && x == 38) || (y == 50 && x == 39) || (y == 51 && x == 39) || (y == 54 && x == 39) || (y == 51 && x == 40) || (y == 51 && x == 42) || (y == 52 && x == 43) || (y == 52 && x == 44) || (y == 53 && x == 44) || (y == 53 && x == 45) || (y == 53 && x == 46) || (y == 55 && x == 46) || (y == 53 && x == 47) || (y == 55 && x == 47) || (y == 53 && x == 48) || (y == 55 && x == 48) || (y == 51 && x == 53) || (y == 52 && x == 53) || (y == 53 && x == 53) || (y == 52 && x == 54) || (y == 51 && x == 55) || (y == 51 && x == 56) || (y == 51 && x == 57) || (y == 50 && x == 58) || (y == 48 && x == 62) || (y == 44 && x == 63) || (y == 47 && x == 63) || (y == 48 && x == 63) || (y == 44 && x == 64) || (y == 46 && x == 64) || (y == 47 && x == 64) || (y == 49 && x == 64) || (y == 50 && x == 64) || (y == 46 && x == 65) || (y == 44 && x == 67) || (y == 45 && x == 67) || (y == 48 && x == 67) || (y == 44 && x == 68) || (y == 47 && x == 68) || (y == 48 && x == 68) || (y == 47 && x == 69) || (y == 47 && x == 70)) oled_data <= 16'h99ce;
        else if ((y == 29 && x == 37)) oled_data <= 16'h2a2c;
        else if ((y == 24 && x == 35)) oled_data <= 16'hd0e1;
        else if ((y == 43 && x == 65) || (y == 41 && x == 71)) oled_data <= 16'ha1ee;
        else if ((y == 42 && x == 36) || (y == 26 && x == 37) || (y == 41 && x == 37) || (y == 40 && x == 54) || (y == 32 && x == 66)) oled_data <= 16'hf880;
        else if ((y == 38 && x == 63)) oled_data <= 16'h490c;
        else if ((y == 38 && x == 69)) oled_data <= 16'h40cf;
        else if ((y == 38 && x == 54)) oled_data <= 16'hc026;
        else if ((y == 37 && x == 58)) oled_data <= 16'h706c;
        else if ((y == 35 && x == 62) || (y == 39 && x == 62)) oled_data <= 16'h414c;
        else if ((y == 47 && x == 41) || (y == 48 && x == 41)) oled_data <= 16'hff74;
        else if ((y == 27 && x == 42)) oled_data <= 16'h226d;
        else if ((y == 41 && x == 31) || (y == 42 && x == 68)) oled_data <= 16'h380b;
        else if ((y == 32 && x == 65)) oled_data <= 16'hf0a0;
        else if ((y == 47 && x == 30)) oled_data <= 16'h79ec;
        else if ((y == 43 && x == 50)) oled_data <= 16'hffba;
        else if ((y == 44 && x == 58)) oled_data <= 16'h5173;
        else if ((y == 25 && x == 30)) oled_data <= 16'h38d2;
        else if ((y == 39 && x == 35)) oled_data <= 16'h263d;
        else if ((y == 22 && x == 35) || (y == 24 && x == 66)) oled_data <= 16'h4076;
        else if ((y == 53 && x == 43) || (y == 53 && x == 49)) oled_data <= 16'h69ec;
        else if ((y == 45 && x == 27) || (y == 45 && x == 64)) oled_data <= 16'h71ec;
        else if ((y == 46 && x == 22) || (y == 47 && x == 26) || (y == 50 && x == 27) || (y == 47 && x == 29) || (y == 53 && x == 33) || (y == 55 && x == 43) || (y == 55 && x == 49) || (y == 55 && x == 51) || (y == 55 && x == 52) || (y == 49 && x == 60) || (y == 49 && x == 66) || (y == 43 && x == 68) || (y == 45 && x == 68) || (y == 44 && x == 69)) oled_data <= 16'h5a0b;
        else if ((y == 44 && x == 33)) oled_data <= 16'h386b;
        else if ((y == 31 && x == 43) || (y == 24 && x == 49) || (y == 24 && x == 50) || (y == 40 && x == 61)) oled_data <= 16'h902a;
        else if ((y == 45 && x == 46)) oled_data <= 16'hddbd;
        else if ((y == 24 && x == 48)) oled_data <= 16'h31ab;
        else if ((y == 35 && x == 38) || (y == 28 && x == 46) || (y == 26 && x == 47) || (y == 35 && x == 56)) oled_data <= 16'h50ad;
        else if ((y == 39 && x == 45) || (y == 40 && x == 50)) oled_data <= 16'hfde0;
        else if ((y == 18 && x == 43) || (y == 18 && x == 54)) oled_data <= 16'h6016;
        else if ((y == 50 && x == 57)) oled_data <= 16'h508d;
        else if ((y == 38 && x == 61) || (y == 40 && x == 62) || (y == 41 && x == 62)) oled_data <= 16'h784b;
        else if ((y == 24 && x == 46) || (y == 26 && x == 55)) oled_data <= 16'h171f;
        else if ((y == 52 && x == 26) || (y == 53 && x == 27) || (y == 54 && x == 28) || (y == 25 && x == 29) || (y == 23 && x == 30) || (y == 16 && x == 38) || (y == 15 && x == 45) || (y == 18 && x == 47) || (y == 57 && x == 47) || (y == 18 && x == 48) || (y == 57 && x == 48) || (y == 18 && x == 49) || (y == 57 && x == 49) || (y == 18 && x == 50) || (y == 9 && x == 51) || (y == 10 && x == 51) || (y == 15 && x == 51) || (y == 9 && x == 52) || (y == 10 && x == 52) || (y == 15 && x == 52) || (y == 15 && x == 56) || (y == 16 && x == 59) || (y == 54 && x == 64) || (y == 23 && x == 65) || (y == 52 && x == 69) || (y == 31 && x == 73) || (y == 48 && x == 73) || (y == 33 && x == 74) || (y == 46 && x == 74)) oled_data <= 16'h29a7;
        else if ((y == 54 && x == 38) || (y == 51 && x == 60)) oled_data <= 16'h59eb;
        else if ((y == 29 && x == 39)) oled_data <= 16'he8c1;
        else if ((y == 34 && x == 39)) oled_data <= 16'h482c;
        else if ((y == 50 && x == 40)) oled_data <= 16'hbb69;
        else if ((y == 45 && x == 54) || (y == 45 && x == 56)) oled_data <= 16'ha24a;
        else if ((y == 43 && x == 37)) oled_data <= 16'h486e;
        else if ((y == 29 && x == 57)) oled_data <= 16'h29ab;
        else if ((y == 37 && x == 61)) oled_data <= 16'hb1e6;
        else if ((y == 48 && x == 53)) oled_data <= 16'hfe61;
        else if ((y == 49 && x == 50)) oled_data <= 16'hffdc;
        else if ((y == 26 && x == 53)) oled_data <= 16'h606c;
        else if ((y == 38 && x == 48) || (y == 50 && x == 51) || (y == 50 && x == 53)) oled_data <= 16'hfe80;
        else if ((y == 34 && x == 72) || (y == 44 && x == 72)) oled_data <= 16'h2097;
        else if ((y == 35 && x == 28) || (y == 34 && x == 67)) oled_data <= 16'h29c8;
        else if ((y == 44 && x == 34)) oled_data <= 16'h404b;
        else if ((y == 49 && x == 59)) oled_data <= 16'hfada;
        else if ((y == 34 && x == 61) || (y == 35 && x == 61) || (y == 36 && x == 61)) oled_data <= 16'h50ec;
        else if ((y == 33 && x == 66)) oled_data <= 16'h19c9;
        else if ((y == 34 && x == 33) || (y == 35 && x == 33) || (y == 36 && x == 33) || (y == 37 && x == 33) || (y == 38 && x == 33) || (y == 39 && x == 33) || (y == 32 && x == 34) || (y == 37 && x == 34) || (y == 38 && x == 34) || (y == 40 && x == 34) || (y == 41 && x == 34) || (y == 42 && x == 34) || (y == 34 && x == 35) || (y == 35 && x == 35) || (y == 36 && x == 35) || (y == 37 && x == 35) || (y == 40 && x == 35) || (y == 41 && x == 35) || (y == 42 && x == 35) || (y == 44 && x == 35) || (y == 33 && x == 36) || (y == 35 && x == 36) || (y == 44 && x == 36) || (y == 46 && x == 36) || (y == 34 && x == 37) || (y == 43 && x == 38) || (y == 33 && x == 40) || (y == 34 && x == 40) || (y == 34 && x == 41) || (y == 28 && x == 42) || (y == 29 && x == 42) || (y == 30 && x == 42) || (y == 31 && x == 42) || (y == 32 && x == 42) || (y == 27 && x == 43) || (y == 28 && x == 43) || (y == 30 && x == 43) || (y == 27 && x == 44) || (y == 26 && x == 45) || (y == 25 && x == 46) || (y == 27 && x == 46) || (y == 25 && x == 47) || (y == 27 && x == 47) || (y == 23 && x == 48) || (y == 26 && x == 48) || (y == 23 && x == 49) || (y == 23 && x == 50) || (y == 25 && x == 50) || (y == 24 && x == 51) || (y == 25 && x == 51) || (y == 25 && x == 52) || (y == 26 && x == 52) || (y == 28 && x == 53) || (y == 29 && x == 54) || (y == 30 && x == 54) || (y == 31 && x == 54) || (y == 27 && x == 55) || (y == 32 && x == 55) || (y == 33 && x == 55) || (y == 35 && x == 55) || (y == 36 && x == 55) || (y == 28 && x == 56) || (y == 49 && x == 56) || (y == 37 && x == 57) || (y == 38 && x == 57) || (y == 49 && x == 57) || (y == 34 && x == 58) || (y == 35 && x == 58) || (y == 36 && x == 58) || (y == 38 && x == 58) || (y == 45 && x == 58) || (y == 46 && x == 58) || (y == 48 && x == 58) || (y == 33 && x == 59) || (y == 34 && x == 59) || (y == 35 && x == 59) || (y == 36 && x == 59) || (y == 37 && x == 59) || (y == 45 && x == 59) || (y == 46 && x == 59) || (y == 31 && x == 60) || (y == 33 && x == 60) || (y == 34 && x == 60) || (y == 35 && x == 60) || (y == 36 && x == 60) || (y == 37 && x == 60) || (y == 44 && x == 60) || (y == 45 && x == 60) || (y == 31 && x == 61) || (y == 32 && x == 61) || (y == 33 && x == 61) || (y == 44 && x == 61) || (y == 45 && x == 61) || (y == 32 && x == 62) || (y == 33 && x == 62) || (y == 34 && x == 62) || (y == 42 && x == 62) || (y == 39 && x == 63) || (y == 40 && x == 63) || (y == 41 && x == 63)) oled_data <= 16'h58ad;
        else if ((y == 33 && x == 41)) oled_data <= 16'h802b;
        else if ((y == 39 && x == 34)) oled_data <= 16'hb9d;
        else if ((y == 45 && x == 43)) oled_data <= 16'h4974;
        else if ((y == 27 && x == 61)) oled_data <= 16'hfaa0;
        else if ((y == 30 && x == 57)) oled_data <= 16'h657f;
        else if ((y == 44 && x == 62)) oled_data <= 16'h510f;
        else if ((y == 24 && x == 31)) oled_data <= 16'h4094;
        else if ((y == 25 && x == 57) || (y == 26 && x == 57) || (y == 27 && x == 57)) oled_data <= 16'h173f;
        else if ((y == 44 && x == 29) || (y == 51 && x == 33)) oled_data <= 16'h31cb;
        else if ((y == 34 && x == 55)) oled_data <= 16'h586c;
        else if ((y == 30 && x == 40)) oled_data <= 16'h9167;
        else if ((y == 45 && x == 47)) oled_data <= 16'hdd9d;
        else if ((y == 52 && x == 48)) oled_data <= 16'hfe1d;
        else if ((y == 51 && x == 37) || (y == 54 && x == 48) || (y == 54 && x == 49) || (y == 51 && x == 58) || (y == 51 && x == 63)) oled_data <= 16'h91cd;
        else if ((y == 52 && x == 45)) oled_data <= 16'hddb9;
        else if ((y == 44 && x == 37) || (y == 49 && x == 38) || (y == 35 && x == 44) || (y == 39 && x == 44) || (y == 34 && x == 45) || (y == 41 && x == 45) || (y == 33 && x == 47) || (y == 33 && x == 48) || (y == 45 && x == 55) || (y == 43 && x == 57) || (y == 47 && x == 57)) oled_data <= 16'hfb20;
        else if ((y == 45 && x == 28)) oled_data <= 16'h61cc;
        else if ((y == 47 && x == 32) || (y == 45 && x == 33) || (y == 47 && x == 33) || (y == 49 && x == 33) || (y == 47 && x == 34) || (y == 47 && x == 35) || (y == 50 && x == 42) || (y == 51 && x == 43) || (y == 51 && x == 46) || (y == 52 && x == 46) || (y == 52 && x == 47) || (y == 52 && x == 49) || (y == 51 && x == 51) || (y == 52 && x == 51) || (y == 53 && x == 51) || (y == 50 && x == 52) || (y == 51 && x == 52) || (y == 48 && x == 60) || (y == 46 && x == 61) || (y == 50 && x == 62)) oled_data <= 16'hfab8;
        else if ((y == 35 && x == 51)) oled_data <= 16'hd044;
        else if ((y == 33 && x == 37)) oled_data <= 16'h175f;
        else if ((y == 37 && x == 26) || (y == 39 && x == 26) || (y == 36 && x == 27) || (y == 37 && x == 27) || (y == 38 && x == 27) || (y == 39 && x == 27) || (y == 40 && x == 27) || (y == 41 && x == 27) || (y == 36 && x == 28) || (y == 39 && x == 28) || (y == 40 && x == 28) || (y == 35 && x == 29) || (y == 40 && x == 29) || (y == 41 && x == 29) || (y == 42 && x == 29) || (y == 35 && x == 30) || (y == 41 && x == 30) || (y == 42 && x == 30) || (y == 43 && x == 30) || (y == 42 && x == 31) || (y == 43 && x == 31) || (y == 42 && x == 32) || (y == 42 && x == 33) || (y == 43 && x == 33) || (y == 43 && x == 34) || (y == 43 && x == 35) || (y == 43 && x == 36) || (y == 43 && x == 60) || (y == 43 && x == 61) || (y == 43 && x == 62) || (y == 42 && x == 63) || (y == 43 && x == 63) || (y == 42 && x == 64) || (y == 43 && x == 64) || (y == 41 && x == 65) || (y == 42 && x == 65) || (y == 40 && x == 66) || (y == 41 && x == 66) || (y == 42 && x == 66) || (y == 43 && x == 66) || (y == 40 && x == 67) || (y == 41 && x == 67) || (y == 42 && x == 67) || (y == 43 && x == 67) || (y == 40 && x == 68) || (y == 41 && x == 68) || (y == 35 && x == 69) || (y == 39 && x == 69) || (y == 40 && x == 69) || (y == 41 && x == 69) || (y == 43 && x == 69) || (y == 36 && x == 70) || (y == 37 && x == 70) || (y == 38 && x == 70) || (y == 39 && x == 70) || (y == 40 && x == 70) || (y == 42 && x == 70) || (y == 37 && x == 71) || (y == 38 && x == 71) || (y == 39 && x == 71) || (y == 40 && x == 71)) oled_data <= 16'h382b;
        else if ((y == 53 && x == 37)) oled_data <= 16'h89cd;
        else if ((y == 46 && x == 44) || (y == 48 && x == 52)) oled_data <= 16'hffb8;
        else if ((y == 41 && x == 51)) oled_data <= 16'hfea0;
        else if ((y == 41 && x == 38) || (y == 46 && x == 39) || (y == 41 && x == 55)) oled_data <= 16'hfb40;
        else if ((y == 33 && x == 26) || (y == 22 && x == 34) || (y == 24 && x == 65) || (y == 27 && x == 68) || (y == 29 && x == 70)) oled_data <= 16'h481b;
        else if ((y == 33 && x == 51) || (y == 34 && x == 51)) oled_data <= 16'hfa00;
        else if ((y == 25 && x == 62) || (y == 28 && x == 62)) oled_data <= 16'h60e9;
        else if ((y == 31 && x == 29) || (y == 29 && x == 61) || (y == 31 && x == 63)) oled_data <= 16'h29ca;
        else if ((y == 23 && x == 34) || (y == 25 && x == 37) || (y == 42 && x == 38) || (y == 36 && x == 40) || (y == 28 && x == 44) || (y == 26 && x == 49) || (y == 26 && x == 50) || (y == 26 && x == 51) || (y == 36 && x == 53) || (y == 33 && x == 58) || (y == 35 && x == 63)) oled_data <= 16'ha809;
        else if ((y == 20 && x == 37)) oled_data <= 16'h29e6;
        else if ((y == 33 && x == 71)) oled_data <= 16'h318a;
        else if ((y == 45 && x == 45)) oled_data <= 16'hbb3a;
        else if ((y == 19 && x == 40) || (y == 20 && x == 59)) oled_data <= 16'h6816;
        else if ((y == 48 && x == 57)) oled_data <= 16'h41f;
        else if ((y == 37 && x == 42) || (y == 42 && x == 44)) oled_data <= 16'hfae0;
        else if ((y == 37 && x == 30)) oled_data <= 16'h39ae;
        else if ((y == 31 && x == 27)) oled_data <= 16'h392e;
        else if ((y == 44 && x == 26)) oled_data <= 16'h39a9;
        else if ((y == 38 && x == 72)) oled_data <= 16'h30aa;
        else if ((y == 36 && x == 29) || (y == 37 && x == 29) || (y == 36 && x == 30) || (y == 35 && x == 31) || (y == 35 && x == 32) || (y == 35 && x == 34) || (y == 44 && x == 38) || (y == 44 && x == 39) || (y == 45 && x == 40) || (y == 45 && x == 41) || (y == 45 && x == 42) || (y == 44 && x == 57) || (y == 35 && x == 64) || (y == 35 && x == 65) || (y == 35 && x == 66) || (y == 35 && x == 67) || (y == 36 && x == 67) || (y == 36 && x == 68) || (y == 37 && x == 68)) oled_data <= 16'h5194;
        else if ((y == 30 && x == 39)) oled_data <= 16'h70aa;
        else if ((y == 48 && x == 23) || (y == 27 && x == 27) || (y == 56 && x == 42) || (y == 55 && x == 61) || (y == 27 && x == 70)) oled_data <= 16'h21a6;
        else if ((y == 29 && x == 28)) oled_data <= 16'h4057;
        else if ((y == 41 && x == 26)) oled_data <= 16'h29e7;
        else if ((y == 48 && x == 37) || (y == 51 && x == 54)) oled_data <= 16'h91af;
        else if ((y == 21 && x == 62) || (y == 22 && x == 62)) oled_data <= 16'h38f0;
        else if ((y == 54 && x == 63)) oled_data <= 16'h31c7;
        else if ((y == 37 && x == 69)) oled_data <= 16'h51b5;
        else if ((y == 32 && x == 40)) oled_data <= 16'h58ee;
        else if ((y == 40 && x == 33) || (y == 36 && x == 34) || (y == 33 && x == 39) || (y == 26 && x == 46) || (y == 27 && x == 54) || (y == 33 && x == 56) || (y == 34 && x == 56) || (y == 50 && x == 56) || (y == 32 && x == 59)) oled_data <= 16'h588d;
        else if ((y == 32 && x == 67)) oled_data <= 16'h9809;
        else if ((y == 53 && x == 62) || (y == 53 && x == 65) || (y == 53 && x == 66)) oled_data <= 16'h39c9;
        else if ((y == 26 && x == 42)) oled_data <= 16'h16df;
        else if ((y == 33 && x == 72)) oled_data <= 16'h2098;
        else if ((y == 42 && x == 37)) oled_data <= 16'hfb60;
        else if ((y == 32 && x == 54) || (y == 33 && x == 54)) oled_data <= 16'h9808;
        else if ((y == 24 && x == 37)) oled_data <= 16'h31aa;
        else if ((y == 33 && x == 33)) oled_data <= 16'h608d;
        else if ((y == 18 && x == 51)) oled_data <= 16'h40ed;
        else if ((y == 40 && x == 52)) oled_data <= 16'hfbe0;
        else if ((y == 51 && x == 61)) oled_data <= 16'hb1f0;
        else if ((y == 45 && x == 36) || (y == 23 && x == 51)) oled_data <= 16'h412c;
        else if ((y == 27 && x == 38)) oled_data <= 16'h19ec;
        else if ((y == 44 && x == 40)) oled_data <= 16'h81ee;
        else if ((y == 29 && x == 38) || (y == 34 && x == 66)) oled_data <= 16'h29eb;
        else if ((y == 32 && x == 26) || (y == 30 && x == 27) || (y == 28 && x == 28) || (y == 27 && x == 29) || (y == 26 && x == 30) || (y == 24 && x == 32) || (y == 23 && x == 33) || (y == 21 && x == 36) || (y == 22 && x == 63) || (y == 23 && x == 64) || (y == 25 && x == 67) || (y == 26 && x == 67) || (y == 28 && x == 69) || (y == 30 && x == 70) || (y == 32 && x == 71)) oled_data <= 16'h481a;
        else if ((y == 46 && x == 45) || (y == 50 && x == 50) || (y == 48 && x == 55) || (y == 33 && x == 65)) oled_data <= 16'hfe40;
        else if ((y == 45 && x == 52)) oled_data <= 16'hdd7d;
        else if ((y == 36 && x == 26) || (y == 38 && x == 26) || (y == 40 && x == 26) || (y == 37 && x == 28) || (y == 38 && x == 28) || (y == 41 && x == 28) || (y == 36 && x == 69) || (y == 42 && x == 69) || (y == 41 && x == 70) || (y == 36 && x == 71)) oled_data <= 16'h384b;
        else if ((y == 25 && x == 53) || (y == 35 && x == 54)) oled_data <= 16'h3df;
        else if ((y == 26 && x == 54)) oled_data <= 16'h177f;
        else if ((y == 30 && x == 59)) oled_data <= 16'h592a;
        else if ((y == 30 && x == 44)) oled_data <= 16'hb8a5;
        else if ((y == 34 && x == 22) || (y == 35 && x == 22) || (y == 36 && x == 22) || (y == 37 && x == 22) || (y == 38 && x == 22) || (y == 39 && x == 22) || (y == 40 && x == 22) || (y == 41 && x == 22) || (y == 42 && x == 22) || (y == 43 && x == 22) || (y == 44 && x == 22) || (y == 45 && x == 22) || (y == 32 && x == 23) || (y == 33 && x == 23) || (y == 34 && x == 23) || (y == 35 && x == 23) || (y == 36 && x == 23) || (y == 37 && x == 23) || (y == 38 && x == 23) || (y == 39 && x == 23) || (y == 40 && x == 23) || (y == 41 && x == 23) || (y == 42 && x == 23) || (y == 43 && x == 23) || (y == 44 && x == 23) || (y == 45 && x == 23) || (y == 47 && x == 23) || (y == 31 && x == 24) || (y == 32 && x == 24) || (y == 33 && x == 24) || (y == 34 && x == 24) || (y == 35 && x == 24) || (y == 36 && x == 24) || (y == 37 && x == 24) || (y == 38 && x == 24) || (y == 39 && x == 24) || (y == 40 && x == 24) || (y == 41 && x == 24) || (y == 42 && x == 24) || (y == 43 && x == 24) || (y == 44 && x == 24) || (y == 45 && x == 24) || (y == 46 && x == 24) || (y == 49 && x == 24) || (y == 30 && x == 25) || (y == 31 && x == 25) || (y == 32 && x == 25) || (y == 38 && x == 25) || (y == 39 && x == 25) || (y == 40 && x == 25) || (y == 41 && x == 25) || (y == 42 && x == 25) || (y == 43 && x == 25) || (y == 46 && x == 25) || (y == 50 && x == 25) || (y == 29 && x == 26) || (y == 30 && x == 26) || (y == 34 && x == 26) || (y == 35 && x == 26) || (y == 42 && x == 26) || (y == 43 && x == 26) || (y == 50 && x == 26) || (y == 51 && x == 26) || (y == 28 && x == 27) || (y == 32 && x == 27) || (y == 33 && x == 27) || (y == 34 && x == 27) || (y == 35 && x == 27) || (y == 51 && x == 27) || (y == 52 && x == 27) || (y == 27 && x == 28) || (y == 30 && x == 28) || (y == 31 && x == 28) || (y == 32 && x == 28) || (y == 33 && x == 28) || (y == 34 && x == 28) || (y == 51 && x == 28) || (y == 52 && x == 28) || (y == 53 && x == 28) || (y == 26 && x == 29) || (y == 28 && x == 29) || (y == 29 && x == 29) || (y == 30 && x == 29) || (y == 51 && x == 29) || (y == 52 && x == 29) || (y == 53 && x == 29) || (y == 54 && x == 29) || (y == 24 && x == 30) || (y == 27 && x == 30) || (y == 28 && x == 30) || (y == 51 && x == 30) || (y == 52 && x == 30) || (y == 53 && x == 30) || (y == 54 && x == 30) || (y == 55 && x == 30) || (y == 22 && x == 31) || (y == 23 && x == 31) || (y == 26 && x == 31) || (y == 27 && x == 31) || (y == 51 && x == 31) || (y == 52 && x == 31) || (y == 53 && x == 31) || (y == 54 && x == 31) || (y == 55 && x == 31) || (y == 56 && x == 31) || (y == 20 && x == 32) || (y == 21 && x == 32) || (y == 22 && x == 32) || (y == 23 && x == 32) || (y == 25 && x == 32) || (y == 26 && x == 32) || (y == 51 && x == 32) || (y == 52 && x == 32) || (y == 53 && x == 32) || (y == 54 && x == 32) || (y == 55 && x == 32) || (y == 56 && x == 32) || (y == 19 && x == 33) || (y == 20 && x == 33) || (y == 21 && x == 33) || (y == 22 && x == 33) || (y == 24 && x == 33) || (y == 25 && x == 33) || (y == 54 && x == 33) || (y == 55 && x == 33) || (y == 56 && x == 33) || (y == 57 && x == 33) || (y == 18 && x == 34) || (y == 19 && x == 34) || (y == 20 && x == 34) || (y == 21 && x == 34) || (y == 24 && x == 34) || (y == 54 && x == 34) || (y == 55 && x == 34) || (y == 56 && x == 34) || (y == 57 && x == 34) || (y == 18 && x == 35) || (y == 19 && x == 35) || (y == 20 && x == 35) || (y == 21 && x == 35) || (y == 54 && x == 35) || (y == 55 && x == 35) || (y == 56 && x == 35) || (y == 57 && x == 35) || (y == 17 && x == 36) || (y == 18 && x == 36) || (y == 19 && x == 36) || (y == 20 && x == 36) || (y == 22 && x == 36) || (y == 23 && x == 36) || (y == 54 && x == 36) || (y == 55 && x == 36) || (y == 56 && x == 36) || (y == 57 && x == 36) || (y == 17 && x == 37) || (y == 18 && x == 37) || (y == 19 && x == 37) || (y == 21 && x == 37) || (y == 22 && x == 37) || (y == 23 && x == 37) || (y == 54 && x == 37) || (y == 55 && x == 37) || (y == 56 && x == 37) || (y == 57 && x == 37) || (y == 17 && x == 38) || (y == 18 && x == 38) || (y == 19 && x == 38) || (y == 21 && x == 38) || (y == 22 && x == 38) || (y == 23 && x == 38) || (y == 53 && x == 38) || (y == 55 && x == 38) || (y == 56 && x == 38) || (y == 57 && x == 38) || (y == 16 && x == 39) || (y == 17 && x == 39) || (y == 18 && x == 39) || (y == 20 && x == 39) || (y == 21 && x == 39) || (y == 22 && x == 39) || (y == 23 && x == 39) || (y == 53 && x == 39) || (y == 56 && x == 39) || (y == 57 && x == 39) || (y == 16 && x == 40) || (y == 17 && x == 40) || (y == 18 && x == 40) || (y == 20 && x == 40) || (y == 21 && x == 40) || (y == 22 && x == 40) || (y == 23 && x == 40) || (y == 54 && x == 40) || (y == 56 && x == 40) || (y == 16 && x == 41) || (y == 17 && x == 41) || (y == 18 && x == 41) || (y == 20 && x == 41) || (y == 21 && x == 41) || (y == 22 && x == 41) || (y == 54 && x == 41) || (y == 55 && x == 41) || (y == 56 && x == 41) || (y == 16 && x == 42) || (y == 17 && x == 42) || (y == 18 && x == 42) || (y == 20 && x == 42) || (y == 21 && x == 42) || (y == 54 && x == 42) || (y == 55 && x == 42) || (y == 16 && x == 43) || (y == 17 && x == 43) || (y == 19 && x == 43) || (y == 20 && x == 43) || (y == 21 && x == 43) || (y == 54 && x == 43) || (y == 56 && x == 43) || (y == 16 && x == 44) || (y == 17 && x == 44) || (y == 19 && x == 44) || (y == 20 && x == 44) || (y == 21 && x == 44) || (y == 56 && x == 44) || (y == 16 && x == 45) || (y == 17 && x == 45) || (y == 19 && x == 45) || (y == 20 && x == 45) || (y == 21 && x == 45) || (y == 56 && x == 45) || (y == 15 && x == 46) || (y == 16 && x == 46) || (y == 17 && x == 46) || (y == 19 && x == 46) || (y == 20 && x == 46) || (y == 15 && x == 47) || (y == 16 && x == 47) || (y == 17 && x == 47) || (y == 19 && x == 47) || (y == 20 && x == 47) || (y == 15 && x == 48) || (y == 16 && x == 48) || (y == 17 && x == 48) || (y == 19 && x == 48) || (y == 20 && x == 48) || (y == 15 && x == 49) || (y == 16 && x == 49) || (y == 17 && x == 49) || (y == 19 && x == 49) || (y == 20 && x == 49) || (y == 21 && x == 49) || (y == 16 && x == 50) || (y == 17 && x == 50) || (y == 19 && x == 50) || (y == 20 && x == 50) || (y == 21 && x == 50) || (y == 55 && x == 50) || (y == 16 && x == 51) || (y == 17 && x == 51) || (y == 19 && x == 51) || (y == 20 && x == 51) || (y == 21 && x == 51) || (y == 16 && x == 52) || (y == 17 && x == 52) || (y == 19 && x == 52) || (y == 20 && x == 52) || (y == 21 && x == 52) || (y == 15 && x == 53) || (y == 16 && x == 53) || (y == 17 && x == 53) || (y == 19 && x == 53) || (y == 20 && x == 53) || (y == 21 && x == 53) || (y == 22 && x == 53) || (y == 56 && x == 53) || (y == 15 && x == 54) || (y == 16 && x == 54) || (y == 17 && x == 54) || (y == 19 && x == 54) || (y == 20 && x == 54) || (y == 21 && x == 54) || (y == 22 && x == 54) || (y == 23 && x == 54) || (y == 54 && x == 54) || (y == 55 && x == 54) || (y == 56 && x == 54) || (y == 15 && x == 55) || (y == 16 && x == 55) || (y == 17 && x == 55) || (y == 20 && x == 55) || (y == 21 && x == 55) || (y == 22 && x == 55) || (y == 23 && x == 55) || (y == 24 && x == 55) || (y == 54 && x == 55) || (y == 55 && x == 55) || (y == 56 && x == 55) || (y == 16 && x == 56) || (y == 17 && x == 56) || (y == 18 && x == 56) || (y == 20 && x == 56) || (y == 21 && x == 56) || (y == 22 && x == 56) || (y == 23 && x == 56) || (y == 24 && x == 56) || (y == 25 && x == 56) || (y == 54 && x == 56) || (y == 56 && x == 56) || (y == 16 && x == 57) || (y == 17 && x == 57) || (y == 18 && x == 57) || (y == 20 && x == 57) || (y == 21 && x == 57) || (y == 22 && x == 57) || (y == 23 && x == 57) || (y == 24 && x == 57) || (y == 56 && x == 57) || (y == 16 && x == 58) || (y == 17 && x == 58) || (y == 18 && x == 58) || (y == 20 && x == 58) || (y == 21 && x == 58) || (y == 22 && x == 58) || (y == 23 && x == 58) || (y == 24 && x == 58) || (y == 25 && x == 58) || (y == 26 && x == 58) || (y == 56 && x == 58) || (y == 17 && x == 59) || (y == 18 && x == 59) || (y == 19 && x == 59) || (y == 21 && x == 59) || (y == 22 && x == 59) || (y == 23 && x == 59) || (y == 24 && x == 59) || (y == 25 && x == 59) || (y == 26 && x == 59) || (y == 27 && x == 59) || (y == 54 && x == 59) || (y == 17 && x == 60) || (y == 18 && x == 60) || (y == 19 && x == 60) || (y == 21 && x == 60) || (y == 22 && x == 60) || (y == 23 && x == 60) || (y == 24 && x == 60) || (y == 25 && x == 60) || (y == 54 && x == 60) || (y == 18 && x == 61) || (y == 19 && x == 61) || (y == 20 && x == 61) || (y == 22 && x == 61) || (y == 23 && x == 61) || (y == 24 && x == 61) || (y == 19 && x == 62) || (y == 20 && x == 62) || (y == 23 && x == 62) || (y == 24 && x == 62) || (y == 29 && x == 62) || (y == 20 && x == 63) || (y == 21 && x == 63) || (y == 23 && x == 63) || (y == 24 && x == 63) || (y == 25 && x == 63) || (y == 26 && x == 63) || (y == 27 && x == 63) || (y == 28 && x == 63) || (y == 29 && x == 63) || (y == 30 && x == 63) || (y == 53 && x == 63) || (y == 21 && x == 64) || (y == 22 && x == 64) || (y == 24 && x == 64) || (y == 25 && x == 64) || (y == 26 && x == 64) || (y == 27 && x == 64) || (y == 28 && x == 64) || (y == 29 && x == 64) || (y == 30 && x == 64) || (y == 31 && x == 64) || (y == 53 && x == 64) || (y == 22 && x == 65) || (y == 25 && x == 65) || (y == 26 && x == 65) || (y == 27 && x == 65) || (y == 28 && x == 65) || (y == 29 && x == 65) || (y == 30 && x == 65) || (y == 31 && x == 65) || (y == 23 && x == 66) || (y == 25 && x == 66) || (y == 26 && x == 66) || (y == 27 && x == 66) || (y == 28 && x == 66) || (y == 29 && x == 66) || (y == 30 && x == 66) || (y == 31 && x == 66) || (y == 27 && x == 67) || (y == 28 && x == 67) || (y == 29 && x == 67) || (y == 30 && x == 67) || (y == 31 && x == 67) || (y == 33 && x == 67) || (y == 53 && x == 67) || (y == 25 && x == 68) || (y == 28 && x == 68) || (y == 29 && x == 68) || (y == 30 && x == 68) || (y == 31 && x == 68) || (y == 32 && x == 68) || (y == 33 && x == 68) || (y == 34 && x == 68) || (y == 50 && x == 68) || (y == 52 && x == 68) || (y == 26 && x == 69) || (y == 27 && x == 69) || (y == 30 && x == 69) || (y == 31 && x == 69) || (y == 32 && x == 69) || (y == 33 && x == 69) || (y == 34 && x == 69) || (y == 45 && x == 69) || (y == 46 && x == 69) || (y == 50 && x == 69) || (y == 51 && x == 69) || (y == 28 && x == 70) || (y == 31 && x == 70) || (y == 32 && x == 70) || (y == 33 && x == 70) || (y == 34 && x == 70) || (y == 35 && x == 70) || (y == 44 && x == 70) || (y == 45 && x == 70) || (y == 46 && x == 70) || (y == 49 && x == 70) || (y == 50 && x == 70) || (y == 51 && x == 70) || (y == 30 && x == 71) || (y == 34 && x == 71) || (y == 35 && x == 71) || (y == 43 && x == 71) || (y == 44 && x == 71) || (y == 46 && x == 71) || (y == 48 && x == 71) || (y == 49 && x == 71) || (y == 50 && x == 71) || (y == 31 && x == 72) || (y == 32 && x == 72) || (y == 39 && x == 72) || (y == 40 && x == 72) || (y == 45 && x == 72) || (y == 46 && x == 72) || (y == 47 && x == 72) || (y == 48 && x == 72) || (y == 49 && x == 72) || (y == 32 && x == 73) || (y == 33 && x == 73) || (y == 34 && x == 73) || (y == 35 && x == 73) || (y == 36 && x == 73) || (y == 42 && x == 73) || (y == 43 && x == 73) || (y == 44 && x == 73) || (y == 45 && x == 73) || (y == 46 && x == 73) || (y == 47 && x == 73) || (y == 34 && x == 74) || (y == 35 && x == 74) || (y == 36 && x == 74) || (y == 37 && x == 74) || (y == 38 && x == 74) || (y == 39 && x == 74) || (y == 40 && x == 74) || (y == 41 && x == 74) || (y == 42 && x == 74) || (y == 43 && x == 74) || (y == 44 && x == 74) || (y == 45 && x == 74)) oled_data <= 16'h31a8;
        else if ((y == 29 && x == 59)) oled_data <= 16'h19cc;
        else if ((y == 44 && x == 55)) oled_data <= 16'hdac3;
        else if ((y == 31 && x == 40)) oled_data <= 16'hc086;
        else if ((y == 31 && x == 59)) oled_data <= 16'h514a;
        else if ((y == 35 && x == 68)) oled_data <= 16'h382a;
        else if ((y == 53 && x == 52)) oled_data <= 16'hca33;
        else if ((y == 29 && x == 53)) oled_data <= 16'h608c;
        else if ((y == 0 && x == 0) || (y == 1 && x == 0) || (y == 2 && x == 0) || (y == 3 && x == 0) || (y == 4 && x == 0) || (y == 5 && x == 0) || (y == 6 && x == 0) || (y == 7 && x == 0) || (y == 8 && x == 0) || (y == 9 && x == 0) || (y == 10 && x == 0) || (y == 11 && x == 0) || (y == 12 && x == 0) || (y == 13 && x == 0) || (y == 14 && x == 0) || (y == 15 && x == 0) || (y == 16 && x == 0) || (y == 17 && x == 0) || (y == 18 && x == 0) || (y == 19 && x == 0) || (y == 20 && x == 0) || (y == 21 && x == 0) || (y == 22 && x == 0) || (y == 23 && x == 0) || (y == 24 && x == 0) || (y == 25 && x == 0) || (y == 26 && x == 0) || (y == 27 && x == 0) || (y == 28 && x == 0) || (y == 29 && x == 0) || (y == 30 && x == 0) || (y == 31 && x == 0) || (y == 32 && x == 0) || (y == 33 && x == 0) || (y == 34 && x == 0) || (y == 35 && x == 0) || (y == 36 && x == 0) || (y == 37 && x == 0) || (y == 38 && x == 0) || (y == 39 && x == 0) || (y == 40 && x == 0) || (y == 41 && x == 0) || (y == 42 && x == 0) || (y == 43 && x == 0) || (y == 44 && x == 0) || (y == 45 && x == 0) || (y == 46 && x == 0) || (y == 47 && x == 0) || (y == 48 && x == 0) || (y == 49 && x == 0) || (y == 50 && x == 0) || (y == 51 && x == 0) || (y == 52 && x == 0) || (y == 53 && x == 0) || (y == 54 && x == 0) || (y == 55 && x == 0) || (y == 56 && x == 0) || (y == 57 && x == 0) || (y == 58 && x == 0) || (y == 59 && x == 0) || (y == 60 && x == 0) || (y == 61 && x == 0) || (y == 62 && x == 0) || (y == 63 && x == 0) || (y == 0 && x == 1) || (y == 1 && x == 1) || (y == 2 && x == 1) || (y == 3 && x == 1) || (y == 4 && x == 1) || (y == 5 && x == 1) || (y == 6 && x == 1) || (y == 7 && x == 1) || (y == 8 && x == 1) || (y == 9 && x == 1) || (y == 10 && x == 1) || (y == 11 && x == 1) || (y == 12 && x == 1) || (y == 13 && x == 1) || (y == 14 && x == 1) || (y == 15 && x == 1) || (y == 16 && x == 1) || (y == 17 && x == 1) || (y == 18 && x == 1) || (y == 19 && x == 1) || (y == 20 && x == 1) || (y == 21 && x == 1) || (y == 22 && x == 1) || (y == 23 && x == 1) || (y == 24 && x == 1) || (y == 25 && x == 1) || (y == 26 && x == 1) || (y == 27 && x == 1) || (y == 28 && x == 1) || (y == 29 && x == 1) || (y == 30 && x == 1) || (y == 31 && x == 1) || (y == 32 && x == 1) || (y == 33 && x == 1) || (y == 34 && x == 1) || (y == 35 && x == 1) || (y == 36 && x == 1) || (y == 37 && x == 1) || (y == 38 && x == 1) || (y == 39 && x == 1) || (y == 40 && x == 1) || (y == 41 && x == 1) || (y == 42 && x == 1) || (y == 43 && x == 1) || (y == 44 && x == 1) || (y == 45 && x == 1) || (y == 46 && x == 1) || (y == 47 && x == 1) || (y == 48 && x == 1) || (y == 49 && x == 1) || (y == 50 && x == 1) || (y == 51 && x == 1) || (y == 52 && x == 1) || (y == 53 && x == 1) || (y == 54 && x == 1) || (y == 55 && x == 1) || (y == 56 && x == 1) || (y == 57 && x == 1) || (y == 58 && x == 1) || (y == 59 && x == 1) || (y == 60 && x == 1) || (y == 61 && x == 1) || (y == 62 && x == 1) || (y == 63 && x == 1) || (y == 0 && x == 2) || (y == 1 && x == 2) || (y == 2 && x == 2) || (y == 3 && x == 2) || (y == 4 && x == 2) || (y == 5 && x == 2) || (y == 6 && x == 2) || (y == 7 && x == 2) || (y == 8 && x == 2) || (y == 9 && x == 2) || (y == 10 && x == 2) || (y == 11 && x == 2) || (y == 12 && x == 2) || (y == 13 && x == 2) || (y == 14 && x == 2) || (y == 15 && x == 2) || (y == 16 && x == 2) || (y == 17 && x == 2) || (y == 18 && x == 2) || (y == 19 && x == 2) || (y == 20 && x == 2) || (y == 21 && x == 2) || (y == 22 && x == 2) || (y == 23 && x == 2) || (y == 24 && x == 2) || (y == 25 && x == 2) || (y == 26 && x == 2) || (y == 27 && x == 2) || (y == 28 && x == 2) || (y == 29 && x == 2) || (y == 30 && x == 2) || (y == 31 && x == 2) || (y == 32 && x == 2) || (y == 33 && x == 2) || (y == 34 && x == 2) || (y == 35 && x == 2) || (y == 36 && x == 2) || (y == 37 && x == 2) || (y == 38 && x == 2) || (y == 39 && x == 2) || (y == 40 && x == 2) || (y == 41 && x == 2) || (y == 42 && x == 2) || (y == 43 && x == 2) || (y == 44 && x == 2) || (y == 45 && x == 2) || (y == 46 && x == 2) || (y == 47 && x == 2) || (y == 48 && x == 2) || (y == 49 && x == 2) || (y == 50 && x == 2) || (y == 51 && x == 2) || (y == 52 && x == 2) || (y == 53 && x == 2) || (y == 54 && x == 2) || (y == 55 && x == 2) || (y == 56 && x == 2) || (y == 57 && x == 2) || (y == 58 && x == 2) || (y == 59 && x == 2) || (y == 60 && x == 2) || (y == 61 && x == 2) || (y == 62 && x == 2) || (y == 63 && x == 2) || (y == 0 && x == 3) || (y == 1 && x == 3) || (y == 2 && x == 3) || (y == 3 && x == 3) || (y == 4 && x == 3) || (y == 5 && x == 3) || (y == 6 && x == 3) || (y == 7 && x == 3) || (y == 8 && x == 3) || (y == 9 && x == 3) || (y == 10 && x == 3) || (y == 11 && x == 3) || (y == 12 && x == 3) || (y == 13 && x == 3) || (y == 14 && x == 3) || (y == 15 && x == 3) || (y == 16 && x == 3) || (y == 17 && x == 3) || (y == 18 && x == 3) || (y == 19 && x == 3) || (y == 20 && x == 3) || (y == 21 && x == 3) || (y == 22 && x == 3) || (y == 23 && x == 3) || (y == 24 && x == 3) || (y == 25 && x == 3) || (y == 26 && x == 3) || (y == 27 && x == 3) || (y == 28 && x == 3) || (y == 29 && x == 3) || (y == 30 && x == 3) || (y == 31 && x == 3) || (y == 32 && x == 3) || (y == 33 && x == 3) || (y == 34 && x == 3) || (y == 35 && x == 3) || (y == 36 && x == 3) || (y == 37 && x == 3) || (y == 38 && x == 3) || (y == 39 && x == 3) || (y == 40 && x == 3) || (y == 41 && x == 3) || (y == 42 && x == 3) || (y == 43 && x == 3) || (y == 44 && x == 3) || (y == 45 && x == 3) || (y == 46 && x == 3) || (y == 47 && x == 3) || (y == 48 && x == 3) || (y == 49 && x == 3) || (y == 50 && x == 3) || (y == 51 && x == 3) || (y == 52 && x == 3) || (y == 53 && x == 3) || (y == 54 && x == 3) || (y == 55 && x == 3) || (y == 56 && x == 3) || (y == 57 && x == 3) || (y == 58 && x == 3) || (y == 59 && x == 3) || (y == 60 && x == 3) || (y == 61 && x == 3) || (y == 62 && x == 3) || (y == 63 && x == 3) || (y == 0 && x == 4) || (y == 1 && x == 4) || (y == 2 && x == 4) || (y == 3 && x == 4) || (y == 4 && x == 4) || (y == 5 && x == 4) || (y == 6 && x == 4) || (y == 7 && x == 4) || (y == 8 && x == 4) || (y == 9 && x == 4) || (y == 10 && x == 4) || (y == 11 && x == 4) || (y == 12 && x == 4) || (y == 13 && x == 4) || (y == 14 && x == 4) || (y == 15 && x == 4) || (y == 16 && x == 4) || (y == 17 && x == 4) || (y == 18 && x == 4) || (y == 19 && x == 4) || (y == 20 && x == 4) || (y == 21 && x == 4) || (y == 22 && x == 4) || (y == 23 && x == 4) || (y == 24 && x == 4) || (y == 25 && x == 4) || (y == 26 && x == 4) || (y == 27 && x == 4) || (y == 28 && x == 4) || (y == 29 && x == 4) || (y == 30 && x == 4) || (y == 31 && x == 4) || (y == 32 && x == 4) || (y == 33 && x == 4) || (y == 34 && x == 4) || (y == 35 && x == 4) || (y == 36 && x == 4) || (y == 37 && x == 4) || (y == 38 && x == 4) || (y == 39 && x == 4) || (y == 40 && x == 4) || (y == 41 && x == 4) || (y == 42 && x == 4) || (y == 43 && x == 4) || (y == 44 && x == 4) || (y == 45 && x == 4) || (y == 46 && x == 4) || (y == 47 && x == 4) || (y == 48 && x == 4) || (y == 49 && x == 4) || (y == 50 && x == 4) || (y == 51 && x == 4) || (y == 52 && x == 4) || (y == 53 && x == 4) || (y == 54 && x == 4) || (y == 55 && x == 4) || (y == 56 && x == 4) || (y == 57 && x == 4) || (y == 58 && x == 4) || (y == 59 && x == 4) || (y == 60 && x == 4) || (y == 61 && x == 4) || (y == 62 && x == 4) || (y == 63 && x == 4) || (y == 0 && x == 5) || (y == 1 && x == 5) || (y == 2 && x == 5) || (y == 3 && x == 5) || (y == 4 && x == 5) || (y == 5 && x == 5) || (y == 6 && x == 5) || (y == 7 && x == 5) || (y == 8 && x == 5) || (y == 9 && x == 5) || (y == 10 && x == 5) || (y == 11 && x == 5) || (y == 12 && x == 5) || (y == 13 && x == 5) || (y == 14 && x == 5) || (y == 15 && x == 5) || (y == 16 && x == 5) || (y == 17 && x == 5) || (y == 18 && x == 5) || (y == 19 && x == 5) || (y == 20 && x == 5) || (y == 21 && x == 5) || (y == 22 && x == 5) || (y == 23 && x == 5) || (y == 24 && x == 5) || (y == 25 && x == 5) || (y == 26 && x == 5) || (y == 27 && x == 5) || (y == 28 && x == 5) || (y == 29 && x == 5) || (y == 30 && x == 5) || (y == 31 && x == 5) || (y == 32 && x == 5) || (y == 33 && x == 5) || (y == 34 && x == 5) || (y == 35 && x == 5) || (y == 36 && x == 5) || (y == 37 && x == 5) || (y == 38 && x == 5) || (y == 39 && x == 5) || (y == 40 && x == 5) || (y == 41 && x == 5) || (y == 42 && x == 5) || (y == 43 && x == 5) || (y == 44 && x == 5) || (y == 45 && x == 5) || (y == 46 && x == 5) || (y == 47 && x == 5) || (y == 48 && x == 5) || (y == 49 && x == 5) || (y == 50 && x == 5) || (y == 51 && x == 5) || (y == 52 && x == 5) || (y == 53 && x == 5) || (y == 54 && x == 5) || (y == 55 && x == 5) || (y == 56 && x == 5) || (y == 57 && x == 5) || (y == 58 && x == 5) || (y == 59 && x == 5) || (y == 60 && x == 5) || (y == 61 && x == 5) || (y == 62 && x == 5) || (y == 63 && x == 5) || (y == 0 && x == 6) || (y == 1 && x == 6) || (y == 2 && x == 6) || (y == 3 && x == 6) || (y == 4 && x == 6) || (y == 5 && x == 6) || (y == 6 && x == 6) || (y == 7 && x == 6) || (y == 8 && x == 6) || (y == 9 && x == 6) || (y == 10 && x == 6) || (y == 11 && x == 6) || (y == 12 && x == 6) || (y == 13 && x == 6) || (y == 14 && x == 6) || (y == 15 && x == 6) || (y == 16 && x == 6) || (y == 17 && x == 6) || (y == 18 && x == 6) || (y == 19 && x == 6) || (y == 20 && x == 6) || (y == 21 && x == 6) || (y == 22 && x == 6) || (y == 23 && x == 6) || (y == 24 && x == 6) || (y == 25 && x == 6) || (y == 26 && x == 6) || (y == 27 && x == 6) || (y == 28 && x == 6) || (y == 29 && x == 6) || (y == 30 && x == 6) || (y == 31 && x == 6) || (y == 32 && x == 6) || (y == 33 && x == 6) || (y == 34 && x == 6) || (y == 35 && x == 6) || (y == 36 && x == 6) || (y == 37 && x == 6) || (y == 38 && x == 6) || (y == 39 && x == 6) || (y == 40 && x == 6) || (y == 41 && x == 6) || (y == 42 && x == 6) || (y == 43 && x == 6) || (y == 44 && x == 6) || (y == 45 && x == 6) || (y == 46 && x == 6) || (y == 47 && x == 6) || (y == 48 && x == 6) || (y == 49 && x == 6) || (y == 50 && x == 6) || (y == 51 && x == 6) || (y == 52 && x == 6) || (y == 53 && x == 6) || (y == 54 && x == 6) || (y == 55 && x == 6) || (y == 56 && x == 6) || (y == 57 && x == 6) || (y == 58 && x == 6) || (y == 59 && x == 6) || (y == 60 && x == 6) || (y == 61 && x == 6) || (y == 62 && x == 6) || (y == 63 && x == 6) || (y == 0 && x == 7) || (y == 1 && x == 7) || (y == 2 && x == 7) || (y == 3 && x == 7) || (y == 4 && x == 7) || (y == 5 && x == 7) || (y == 6 && x == 7) || (y == 7 && x == 7) || (y == 8 && x == 7) || (y == 9 && x == 7) || (y == 10 && x == 7) || (y == 11 && x == 7) || (y == 12 && x == 7) || (y == 13 && x == 7) || (y == 14 && x == 7) || (y == 15 && x == 7) || (y == 16 && x == 7) || (y == 17 && x == 7) || (y == 18 && x == 7) || (y == 19 && x == 7) || (y == 20 && x == 7) || (y == 21 && x == 7) || (y == 22 && x == 7) || (y == 23 && x == 7) || (y == 24 && x == 7) || (y == 25 && x == 7) || (y == 26 && x == 7) || (y == 27 && x == 7) || (y == 28 && x == 7) || (y == 29 && x == 7) || (y == 30 && x == 7) || (y == 31 && x == 7) || (y == 32 && x == 7) || (y == 33 && x == 7) || (y == 34 && x == 7) || (y == 35 && x == 7) || (y == 36 && x == 7) || (y == 37 && x == 7) || (y == 38 && x == 7) || (y == 39 && x == 7) || (y == 40 && x == 7) || (y == 41 && x == 7) || (y == 42 && x == 7) || (y == 43 && x == 7) || (y == 44 && x == 7) || (y == 45 && x == 7) || (y == 46 && x == 7) || (y == 47 && x == 7) || (y == 48 && x == 7) || (y == 49 && x == 7) || (y == 50 && x == 7) || (y == 51 && x == 7) || (y == 52 && x == 7) || (y == 53 && x == 7) || (y == 54 && x == 7) || (y == 55 && x == 7) || (y == 56 && x == 7) || (y == 57 && x == 7) || (y == 58 && x == 7) || (y == 59 && x == 7) || (y == 60 && x == 7) || (y == 61 && x == 7) || (y == 62 && x == 7) || (y == 63 && x == 7) || (y == 0 && x == 8) || (y == 1 && x == 8) || (y == 2 && x == 8) || (y == 3 && x == 8) || (y == 4 && x == 8) || (y == 5 && x == 8) || (y == 6 && x == 8) || (y == 7 && x == 8) || (y == 8 && x == 8) || (y == 9 && x == 8) || (y == 10 && x == 8) || (y == 11 && x == 8) || (y == 12 && x == 8) || (y == 13 && x == 8) || (y == 14 && x == 8) || (y == 15 && x == 8) || (y == 16 && x == 8) || (y == 17 && x == 8) || (y == 18 && x == 8) || (y == 19 && x == 8) || (y == 20 && x == 8) || (y == 21 && x == 8) || (y == 22 && x == 8) || (y == 23 && x == 8) || (y == 24 && x == 8) || (y == 25 && x == 8) || (y == 26 && x == 8) || (y == 27 && x == 8) || (y == 28 && x == 8) || (y == 29 && x == 8) || (y == 30 && x == 8) || (y == 31 && x == 8) || (y == 32 && x == 8) || (y == 33 && x == 8) || (y == 34 && x == 8) || (y == 35 && x == 8) || (y == 36 && x == 8) || (y == 37 && x == 8) || (y == 38 && x == 8) || (y == 39 && x == 8) || (y == 40 && x == 8) || (y == 41 && x == 8) || (y == 42 && x == 8) || (y == 43 && x == 8) || (y == 44 && x == 8) || (y == 45 && x == 8) || (y == 46 && x == 8) || (y == 47 && x == 8) || (y == 48 && x == 8) || (y == 49 && x == 8) || (y == 50 && x == 8) || (y == 51 && x == 8) || (y == 52 && x == 8) || (y == 53 && x == 8) || (y == 54 && x == 8) || (y == 55 && x == 8) || (y == 56 && x == 8) || (y == 57 && x == 8) || (y == 58 && x == 8) || (y == 59 && x == 8) || (y == 60 && x == 8) || (y == 61 && x == 8) || (y == 62 && x == 8) || (y == 63 && x == 8) || (y == 0 && x == 9) || (y == 1 && x == 9) || (y == 2 && x == 9) || (y == 3 && x == 9) || (y == 4 && x == 9) || (y == 5 && x == 9) || (y == 6 && x == 9) || (y == 7 && x == 9) || (y == 8 && x == 9) || (y == 9 && x == 9) || (y == 10 && x == 9) || (y == 11 && x == 9) || (y == 12 && x == 9) || (y == 13 && x == 9) || (y == 14 && x == 9) || (y == 15 && x == 9) || (y == 16 && x == 9) || (y == 17 && x == 9) || (y == 18 && x == 9) || (y == 19 && x == 9) || (y == 20 && x == 9) || (y == 21 && x == 9) || (y == 22 && x == 9) || (y == 23 && x == 9) || (y == 24 && x == 9) || (y == 25 && x == 9) || (y == 26 && x == 9) || (y == 27 && x == 9) || (y == 28 && x == 9) || (y == 29 && x == 9) || (y == 30 && x == 9) || (y == 31 && x == 9) || (y == 32 && x == 9) || (y == 33 && x == 9) || (y == 34 && x == 9) || (y == 35 && x == 9) || (y == 36 && x == 9) || (y == 37 && x == 9) || (y == 38 && x == 9) || (y == 39 && x == 9) || (y == 40 && x == 9) || (y == 41 && x == 9) || (y == 42 && x == 9) || (y == 43 && x == 9) || (y == 44 && x == 9) || (y == 45 && x == 9) || (y == 46 && x == 9) || (y == 47 && x == 9) || (y == 48 && x == 9) || (y == 49 && x == 9) || (y == 50 && x == 9) || (y == 51 && x == 9) || (y == 52 && x == 9) || (y == 53 && x == 9) || (y == 54 && x == 9) || (y == 55 && x == 9) || (y == 56 && x == 9) || (y == 57 && x == 9) || (y == 58 && x == 9) || (y == 59 && x == 9) || (y == 60 && x == 9) || (y == 61 && x == 9) || (y == 62 && x == 9) || (y == 63 && x == 9) || (y == 0 && x == 10) || (y == 1 && x == 10) || (y == 2 && x == 10) || (y == 3 && x == 10) || (y == 4 && x == 10) || (y == 5 && x == 10) || (y == 6 && x == 10) || (y == 7 && x == 10) || (y == 8 && x == 10) || (y == 9 && x == 10) || (y == 10 && x == 10) || (y == 11 && x == 10) || (y == 12 && x == 10) || (y == 13 && x == 10) || (y == 14 && x == 10) || (y == 15 && x == 10) || (y == 16 && x == 10) || (y == 17 && x == 10) || (y == 18 && x == 10) || (y == 19 && x == 10) || (y == 20 && x == 10) || (y == 21 && x == 10) || (y == 22 && x == 10) || (y == 23 && x == 10) || (y == 24 && x == 10) || (y == 25 && x == 10) || (y == 26 && x == 10) || (y == 27 && x == 10) || (y == 28 && x == 10) || (y == 29 && x == 10) || (y == 30 && x == 10) || (y == 31 && x == 10) || (y == 32 && x == 10) || (y == 33 && x == 10) || (y == 34 && x == 10) || (y == 35 && x == 10) || (y == 36 && x == 10) || (y == 37 && x == 10) || (y == 38 && x == 10) || (y == 39 && x == 10) || (y == 40 && x == 10) || (y == 41 && x == 10) || (y == 42 && x == 10) || (y == 43 && x == 10) || (y == 44 && x == 10) || (y == 45 && x == 10) || (y == 46 && x == 10) || (y == 47 && x == 10) || (y == 48 && x == 10) || (y == 49 && x == 10) || (y == 50 && x == 10) || (y == 51 && x == 10) || (y == 52 && x == 10) || (y == 53 && x == 10) || (y == 54 && x == 10) || (y == 55 && x == 10) || (y == 56 && x == 10) || (y == 57 && x == 10) || (y == 58 && x == 10) || (y == 59 && x == 10) || (y == 60 && x == 10) || (y == 61 && x == 10) || (y == 62 && x == 10) || (y == 63 && x == 10) || (y == 0 && x == 11) || (y == 1 && x == 11) || (y == 2 && x == 11) || (y == 3 && x == 11) || (y == 4 && x == 11) || (y == 5 && x == 11) || (y == 6 && x == 11) || (y == 7 && x == 11) || (y == 8 && x == 11) || (y == 9 && x == 11) || (y == 10 && x == 11) || (y == 11 && x == 11) || (y == 12 && x == 11) || (y == 13 && x == 11) || (y == 14 && x == 11) || (y == 15 && x == 11) || (y == 16 && x == 11) || (y == 17 && x == 11) || (y == 18 && x == 11) || (y == 19 && x == 11) || (y == 20 && x == 11) || (y == 21 && x == 11) || (y == 22 && x == 11) || (y == 23 && x == 11) || (y == 24 && x == 11) || (y == 25 && x == 11) || (y == 26 && x == 11) || (y == 27 && x == 11) || (y == 28 && x == 11) || (y == 29 && x == 11) || (y == 30 && x == 11) || (y == 31 && x == 11) || (y == 32 && x == 11) || (y == 33 && x == 11) || (y == 34 && x == 11) || (y == 35 && x == 11) || (y == 36 && x == 11) || (y == 37 && x == 11) || (y == 38 && x == 11) || (y == 39 && x == 11) || (y == 40 && x == 11) || (y == 41 && x == 11) || (y == 42 && x == 11) || (y == 43 && x == 11) || (y == 44 && x == 11) || (y == 45 && x == 11) || (y == 46 && x == 11) || (y == 47 && x == 11) || (y == 48 && x == 11) || (y == 49 && x == 11) || (y == 50 && x == 11) || (y == 51 && x == 11) || (y == 52 && x == 11) || (y == 53 && x == 11) || (y == 54 && x == 11) || (y == 55 && x == 11) || (y == 56 && x == 11) || (y == 57 && x == 11) || (y == 58 && x == 11) || (y == 59 && x == 11) || (y == 60 && x == 11) || (y == 61 && x == 11) || (y == 62 && x == 11) || (y == 63 && x == 11) || (y == 0 && x == 12) || (y == 1 && x == 12) || (y == 2 && x == 12) || (y == 3 && x == 12) || (y == 4 && x == 12) || (y == 5 && x == 12) || (y == 6 && x == 12) || (y == 7 && x == 12) || (y == 8 && x == 12) || (y == 9 && x == 12) || (y == 10 && x == 12) || (y == 11 && x == 12) || (y == 12 && x == 12) || (y == 13 && x == 12) || (y == 14 && x == 12) || (y == 15 && x == 12) || (y == 16 && x == 12) || (y == 17 && x == 12) || (y == 18 && x == 12) || (y == 19 && x == 12) || (y == 20 && x == 12) || (y == 21 && x == 12) || (y == 22 && x == 12) || (y == 23 && x == 12) || (y == 24 && x == 12) || (y == 25 && x == 12) || (y == 26 && x == 12) || (y == 27 && x == 12) || (y == 28 && x == 12) || (y == 29 && x == 12) || (y == 30 && x == 12) || (y == 31 && x == 12) || (y == 32 && x == 12) || (y == 33 && x == 12) || (y == 34 && x == 12) || (y == 35 && x == 12) || (y == 36 && x == 12) || (y == 37 && x == 12) || (y == 38 && x == 12) || (y == 39 && x == 12) || (y == 40 && x == 12) || (y == 41 && x == 12) || (y == 42 && x == 12) || (y == 43 && x == 12) || (y == 44 && x == 12) || (y == 45 && x == 12) || (y == 46 && x == 12) || (y == 47 && x == 12) || (y == 48 && x == 12) || (y == 49 && x == 12) || (y == 50 && x == 12) || (y == 51 && x == 12) || (y == 52 && x == 12) || (y == 53 && x == 12) || (y == 54 && x == 12) || (y == 55 && x == 12) || (y == 56 && x == 12) || (y == 57 && x == 12) || (y == 58 && x == 12) || (y == 59 && x == 12) || (y == 60 && x == 12) || (y == 61 && x == 12) || (y == 62 && x == 12) || (y == 63 && x == 12) || (y == 0 && x == 13) || (y == 1 && x == 13) || (y == 2 && x == 13) || (y == 3 && x == 13) || (y == 4 && x == 13) || (y == 5 && x == 13) || (y == 6 && x == 13) || (y == 7 && x == 13) || (y == 8 && x == 13) || (y == 9 && x == 13) || (y == 10 && x == 13) || (y == 11 && x == 13) || (y == 12 && x == 13) || (y == 13 && x == 13) || (y == 14 && x == 13) || (y == 15 && x == 13) || (y == 16 && x == 13) || (y == 17 && x == 13) || (y == 18 && x == 13) || (y == 19 && x == 13) || (y == 20 && x == 13) || (y == 21 && x == 13) || (y == 22 && x == 13) || (y == 23 && x == 13) || (y == 24 && x == 13) || (y == 25 && x == 13) || (y == 26 && x == 13) || (y == 27 && x == 13) || (y == 28 && x == 13) || (y == 29 && x == 13) || (y == 30 && x == 13) || (y == 31 && x == 13) || (y == 32 && x == 13) || (y == 33 && x == 13) || (y == 34 && x == 13) || (y == 35 && x == 13) || (y == 36 && x == 13) || (y == 37 && x == 13) || (y == 38 && x == 13) || (y == 39 && x == 13) || (y == 40 && x == 13) || (y == 41 && x == 13) || (y == 42 && x == 13) || (y == 43 && x == 13) || (y == 44 && x == 13) || (y == 45 && x == 13) || (y == 46 && x == 13) || (y == 47 && x == 13) || (y == 48 && x == 13) || (y == 49 && x == 13) || (y == 50 && x == 13) || (y == 51 && x == 13) || (y == 52 && x == 13) || (y == 53 && x == 13) || (y == 54 && x == 13) || (y == 55 && x == 13) || (y == 56 && x == 13) || (y == 57 && x == 13) || (y == 58 && x == 13) || (y == 59 && x == 13) || (y == 60 && x == 13) || (y == 61 && x == 13) || (y == 62 && x == 13) || (y == 63 && x == 13) || (y == 0 && x == 14) || (y == 1 && x == 14) || (y == 2 && x == 14) || (y == 3 && x == 14) || (y == 4 && x == 14) || (y == 5 && x == 14) || (y == 6 && x == 14) || (y == 7 && x == 14) || (y == 8 && x == 14) || (y == 9 && x == 14) || (y == 10 && x == 14) || (y == 11 && x == 14) || (y == 12 && x == 14) || (y == 13 && x == 14) || (y == 14 && x == 14) || (y == 15 && x == 14) || (y == 16 && x == 14) || (y == 17 && x == 14) || (y == 18 && x == 14) || (y == 19 && x == 14) || (y == 20 && x == 14) || (y == 21 && x == 14) || (y == 22 && x == 14) || (y == 23 && x == 14) || (y == 24 && x == 14) || (y == 25 && x == 14) || (y == 26 && x == 14) || (y == 27 && x == 14) || (y == 28 && x == 14) || (y == 29 && x == 14) || (y == 30 && x == 14) || (y == 31 && x == 14) || (y == 32 && x == 14) || (y == 33 && x == 14) || (y == 34 && x == 14) || (y == 35 && x == 14) || (y == 36 && x == 14) || (y == 37 && x == 14) || (y == 38 && x == 14) || (y == 39 && x == 14) || (y == 40 && x == 14) || (y == 41 && x == 14) || (y == 42 && x == 14) || (y == 43 && x == 14) || (y == 44 && x == 14) || (y == 45 && x == 14) || (y == 46 && x == 14) || (y == 47 && x == 14) || (y == 48 && x == 14) || (y == 49 && x == 14) || (y == 50 && x == 14) || (y == 51 && x == 14) || (y == 52 && x == 14) || (y == 53 && x == 14) || (y == 54 && x == 14) || (y == 55 && x == 14) || (y == 56 && x == 14) || (y == 57 && x == 14) || (y == 58 && x == 14) || (y == 59 && x == 14) || (y == 60 && x == 14) || (y == 61 && x == 14) || (y == 62 && x == 14) || (y == 63 && x == 14) || (y == 0 && x == 15) || (y == 1 && x == 15) || (y == 2 && x == 15) || (y == 3 && x == 15) || (y == 4 && x == 15) || (y == 5 && x == 15) || (y == 6 && x == 15) || (y == 7 && x == 15) || (y == 8 && x == 15) || (y == 9 && x == 15) || (y == 10 && x == 15) || (y == 11 && x == 15) || (y == 12 && x == 15) || (y == 13 && x == 15) || (y == 14 && x == 15) || (y == 15 && x == 15) || (y == 16 && x == 15) || (y == 17 && x == 15) || (y == 18 && x == 15) || (y == 19 && x == 15) || (y == 20 && x == 15) || (y == 21 && x == 15) || (y == 22 && x == 15) || (y == 23 && x == 15) || (y == 24 && x == 15) || (y == 25 && x == 15) || (y == 26 && x == 15) || (y == 27 && x == 15) || (y == 28 && x == 15) || (y == 29 && x == 15) || (y == 30 && x == 15) || (y == 31 && x == 15) || (y == 32 && x == 15) || (y == 33 && x == 15) || (y == 34 && x == 15) || (y == 35 && x == 15) || (y == 36 && x == 15) || (y == 37 && x == 15) || (y == 38 && x == 15) || (y == 39 && x == 15) || (y == 40 && x == 15) || (y == 41 && x == 15) || (y == 42 && x == 15) || (y == 43 && x == 15) || (y == 44 && x == 15) || (y == 45 && x == 15) || (y == 46 && x == 15) || (y == 47 && x == 15) || (y == 48 && x == 15) || (y == 49 && x == 15) || (y == 50 && x == 15) || (y == 51 && x == 15) || (y == 52 && x == 15) || (y == 53 && x == 15) || (y == 54 && x == 15) || (y == 55 && x == 15) || (y == 56 && x == 15) || (y == 57 && x == 15) || (y == 58 && x == 15) || (y == 59 && x == 15) || (y == 60 && x == 15) || (y == 61 && x == 15) || (y == 62 && x == 15) || (y == 63 && x == 15) || (y == 0 && x == 16) || (y == 1 && x == 16) || (y == 2 && x == 16) || (y == 3 && x == 16) || (y == 4 && x == 16) || (y == 5 && x == 16) || (y == 6 && x == 16) || (y == 7 && x == 16) || (y == 8 && x == 16) || (y == 9 && x == 16) || (y == 10 && x == 16) || (y == 11 && x == 16) || (y == 12 && x == 16) || (y == 13 && x == 16) || (y == 14 && x == 16) || (y == 15 && x == 16) || (y == 16 && x == 16) || (y == 17 && x == 16) || (y == 18 && x == 16) || (y == 19 && x == 16) || (y == 20 && x == 16) || (y == 21 && x == 16) || (y == 22 && x == 16) || (y == 23 && x == 16) || (y == 24 && x == 16) || (y == 25 && x == 16) || (y == 26 && x == 16) || (y == 27 && x == 16) || (y == 28 && x == 16) || (y == 29 && x == 16) || (y == 30 && x == 16) || (y == 31 && x == 16) || (y == 32 && x == 16) || (y == 33 && x == 16) || (y == 34 && x == 16) || (y == 35 && x == 16) || (y == 36 && x == 16) || (y == 37 && x == 16) || (y == 38 && x == 16) || (y == 39 && x == 16) || (y == 40 && x == 16) || (y == 41 && x == 16) || (y == 42 && x == 16) || (y == 43 && x == 16) || (y == 44 && x == 16) || (y == 45 && x == 16) || (y == 46 && x == 16) || (y == 47 && x == 16) || (y == 48 && x == 16) || (y == 49 && x == 16) || (y == 50 && x == 16) || (y == 51 && x == 16) || (y == 52 && x == 16) || (y == 53 && x == 16) || (y == 54 && x == 16) || (y == 55 && x == 16) || (y == 56 && x == 16) || (y == 57 && x == 16) || (y == 58 && x == 16) || (y == 59 && x == 16) || (y == 60 && x == 16) || (y == 61 && x == 16) || (y == 62 && x == 16) || (y == 63 && x == 16) || (y == 0 && x == 17) || (y == 1 && x == 17) || (y == 2 && x == 17) || (y == 3 && x == 17) || (y == 4 && x == 17) || (y == 5 && x == 17) || (y == 6 && x == 17) || (y == 7 && x == 17) || (y == 8 && x == 17) || (y == 9 && x == 17) || (y == 10 && x == 17) || (y == 11 && x == 17) || (y == 12 && x == 17) || (y == 13 && x == 17) || (y == 14 && x == 17) || (y == 15 && x == 17) || (y == 16 && x == 17) || (y == 17 && x == 17) || (y == 18 && x == 17) || (y == 19 && x == 17) || (y == 20 && x == 17) || (y == 21 && x == 17) || (y == 22 && x == 17) || (y == 23 && x == 17) || (y == 24 && x == 17) || (y == 25 && x == 17) || (y == 26 && x == 17) || (y == 27 && x == 17) || (y == 28 && x == 17) || (y == 29 && x == 17) || (y == 30 && x == 17) || (y == 31 && x == 17) || (y == 32 && x == 17) || (y == 33 && x == 17) || (y == 34 && x == 17) || (y == 35 && x == 17) || (y == 36 && x == 17) || (y == 37 && x == 17) || (y == 38 && x == 17) || (y == 39 && x == 17) || (y == 40 && x == 17) || (y == 41 && x == 17) || (y == 42 && x == 17) || (y == 43 && x == 17) || (y == 44 && x == 17) || (y == 45 && x == 17) || (y == 46 && x == 17) || (y == 47 && x == 17) || (y == 48 && x == 17) || (y == 49 && x == 17) || (y == 50 && x == 17) || (y == 51 && x == 17) || (y == 52 && x == 17) || (y == 53 && x == 17) || (y == 54 && x == 17) || (y == 55 && x == 17) || (y == 56 && x == 17) || (y == 57 && x == 17) || (y == 58 && x == 17) || (y == 59 && x == 17) || (y == 60 && x == 17) || (y == 61 && x == 17) || (y == 62 && x == 17) || (y == 63 && x == 17) || (y == 0 && x == 18) || (y == 1 && x == 18) || (y == 2 && x == 18) || (y == 3 && x == 18) || (y == 4 && x == 18) || (y == 5 && x == 18) || (y == 6 && x == 18) || (y == 7 && x == 18) || (y == 8 && x == 18) || (y == 9 && x == 18) || (y == 10 && x == 18) || (y == 11 && x == 18) || (y == 12 && x == 18) || (y == 13 && x == 18) || (y == 14 && x == 18) || (y == 15 && x == 18) || (y == 16 && x == 18) || (y == 17 && x == 18) || (y == 18 && x == 18) || (y == 19 && x == 18) || (y == 20 && x == 18) || (y == 21 && x == 18) || (y == 22 && x == 18) || (y == 23 && x == 18) || (y == 24 && x == 18) || (y == 25 && x == 18) || (y == 26 && x == 18) || (y == 27 && x == 18) || (y == 28 && x == 18) || (y == 29 && x == 18) || (y == 30 && x == 18) || (y == 31 && x == 18) || (y == 32 && x == 18) || (y == 33 && x == 18) || (y == 34 && x == 18) || (y == 35 && x == 18) || (y == 36 && x == 18) || (y == 37 && x == 18) || (y == 38 && x == 18) || (y == 39 && x == 18) || (y == 40 && x == 18) || (y == 41 && x == 18) || (y == 42 && x == 18) || (y == 43 && x == 18) || (y == 44 && x == 18) || (y == 45 && x == 18) || (y == 46 && x == 18) || (y == 47 && x == 18) || (y == 48 && x == 18) || (y == 49 && x == 18) || (y == 50 && x == 18) || (y == 51 && x == 18) || (y == 52 && x == 18) || (y == 53 && x == 18) || (y == 54 && x == 18) || (y == 55 && x == 18) || (y == 56 && x == 18) || (y == 57 && x == 18) || (y == 58 && x == 18) || (y == 59 && x == 18) || (y == 60 && x == 18) || (y == 61 && x == 18) || (y == 62 && x == 18) || (y == 63 && x == 18) || (y == 0 && x == 19) || (y == 1 && x == 19) || (y == 2 && x == 19) || (y == 3 && x == 19) || (y == 4 && x == 19) || (y == 5 && x == 19) || (y == 6 && x == 19) || (y == 7 && x == 19) || (y == 8 && x == 19) || (y == 9 && x == 19) || (y == 10 && x == 19) || (y == 11 && x == 19) || (y == 12 && x == 19) || (y == 13 && x == 19) || (y == 14 && x == 19) || (y == 15 && x == 19) || (y == 16 && x == 19) || (y == 17 && x == 19) || (y == 18 && x == 19) || (y == 19 && x == 19) || (y == 20 && x == 19) || (y == 21 && x == 19) || (y == 22 && x == 19) || (y == 23 && x == 19) || (y == 24 && x == 19) || (y == 25 && x == 19) || (y == 26 && x == 19) || (y == 27 && x == 19) || (y == 28 && x == 19) || (y == 29 && x == 19) || (y == 30 && x == 19) || (y == 31 && x == 19) || (y == 32 && x == 19) || (y == 33 && x == 19) || (y == 34 && x == 19) || (y == 35 && x == 19) || (y == 36 && x == 19) || (y == 37 && x == 19) || (y == 38 && x == 19) || (y == 39 && x == 19) || (y == 40 && x == 19) || (y == 41 && x == 19) || (y == 42 && x == 19) || (y == 43 && x == 19) || (y == 44 && x == 19) || (y == 45 && x == 19) || (y == 46 && x == 19) || (y == 47 && x == 19) || (y == 48 && x == 19) || (y == 49 && x == 19) || (y == 50 && x == 19) || (y == 51 && x == 19) || (y == 52 && x == 19) || (y == 53 && x == 19) || (y == 54 && x == 19) || (y == 55 && x == 19) || (y == 56 && x == 19) || (y == 57 && x == 19) || (y == 58 && x == 19) || (y == 59 && x == 19) || (y == 60 && x == 19) || (y == 61 && x == 19) || (y == 62 && x == 19) || (y == 63 && x == 19) || (y == 0 && x == 20) || (y == 1 && x == 20) || (y == 2 && x == 20) || (y == 3 && x == 20) || (y == 4 && x == 20) || (y == 5 && x == 20) || (y == 6 && x == 20) || (y == 7 && x == 20) || (y == 8 && x == 20) || (y == 9 && x == 20) || (y == 10 && x == 20) || (y == 11 && x == 20) || (y == 12 && x == 20) || (y == 13 && x == 20) || (y == 14 && x == 20) || (y == 15 && x == 20) || (y == 16 && x == 20) || (y == 17 && x == 20) || (y == 18 && x == 20) || (y == 19 && x == 20) || (y == 20 && x == 20) || (y == 21 && x == 20) || (y == 22 && x == 20) || (y == 23 && x == 20) || (y == 24 && x == 20) || (y == 25 && x == 20) || (y == 26 && x == 20) || (y == 27 && x == 20) || (y == 28 && x == 20) || (y == 29 && x == 20) || (y == 30 && x == 20) || (y == 31 && x == 20) || (y == 32 && x == 20) || (y == 33 && x == 20) || (y == 34 && x == 20) || (y == 35 && x == 20) || (y == 36 && x == 20) || (y == 37 && x == 20) || (y == 38 && x == 20) || (y == 39 && x == 20) || (y == 40 && x == 20) || (y == 41 && x == 20) || (y == 42 && x == 20) || (y == 43 && x == 20) || (y == 44 && x == 20) || (y == 45 && x == 20) || (y == 46 && x == 20) || (y == 47 && x == 20) || (y == 48 && x == 20) || (y == 49 && x == 20) || (y == 50 && x == 20) || (y == 51 && x == 20) || (y == 52 && x == 20) || (y == 53 && x == 20) || (y == 54 && x == 20) || (y == 55 && x == 20) || (y == 56 && x == 20) || (y == 57 && x == 20) || (y == 58 && x == 20) || (y == 59 && x == 20) || (y == 60 && x == 20) || (y == 61 && x == 20) || (y == 62 && x == 20) || (y == 63 && x == 20) || (y == 0 && x == 21) || (y == 1 && x == 21) || (y == 2 && x == 21) || (y == 3 && x == 21) || (y == 4 && x == 21) || (y == 5 && x == 21) || (y == 6 && x == 21) || (y == 7 && x == 21) || (y == 8 && x == 21) || (y == 9 && x == 21) || (y == 10 && x == 21) || (y == 11 && x == 21) || (y == 12 && x == 21) || (y == 13 && x == 21) || (y == 14 && x == 21) || (y == 15 && x == 21) || (y == 16 && x == 21) || (y == 17 && x == 21) || (y == 18 && x == 21) || (y == 19 && x == 21) || (y == 20 && x == 21) || (y == 21 && x == 21) || (y == 22 && x == 21) || (y == 23 && x == 21) || (y == 24 && x == 21) || (y == 25 && x == 21) || (y == 26 && x == 21) || (y == 27 && x == 21) || (y == 28 && x == 21) || (y == 29 && x == 21) || (y == 30 && x == 21) || (y == 31 && x == 21) || (y == 32 && x == 21) || (y == 33 && x == 21) || (y == 34 && x == 21) || (y == 35 && x == 21) || (y == 36 && x == 21) || (y == 37 && x == 21) || (y == 38 && x == 21) || (y == 39 && x == 21) || (y == 40 && x == 21) || (y == 41 && x == 21) || (y == 42 && x == 21) || (y == 43 && x == 21) || (y == 44 && x == 21) || (y == 45 && x == 21) || (y == 46 && x == 21) || (y == 47 && x == 21) || (y == 48 && x == 21) || (y == 49 && x == 21) || (y == 50 && x == 21) || (y == 51 && x == 21) || (y == 52 && x == 21) || (y == 53 && x == 21) || (y == 54 && x == 21) || (y == 55 && x == 21) || (y == 56 && x == 21) || (y == 57 && x == 21) || (y == 58 && x == 21) || (y == 59 && x == 21) || (y == 60 && x == 21) || (y == 61 && x == 21) || (y == 62 && x == 21) || (y == 63 && x == 21) || (y == 0 && x == 22) || (y == 1 && x == 22) || (y == 2 && x == 22) || (y == 3 && x == 22) || (y == 4 && x == 22) || (y == 5 && x == 22) || (y == 6 && x == 22) || (y == 7 && x == 22) || (y == 8 && x == 22) || (y == 9 && x == 22) || (y == 10 && x == 22) || (y == 11 && x == 22) || (y == 12 && x == 22) || (y == 13 && x == 22) || (y == 14 && x == 22) || (y == 15 && x == 22) || (y == 16 && x == 22) || (y == 17 && x == 22) || (y == 18 && x == 22) || (y == 19 && x == 22) || (y == 20 && x == 22) || (y == 21 && x == 22) || (y == 22 && x == 22) || (y == 23 && x == 22) || (y == 24 && x == 22) || (y == 25 && x == 22) || (y == 26 && x == 22) || (y == 27 && x == 22) || (y == 28 && x == 22) || (y == 29 && x == 22) || (y == 30 && x == 22) || (y == 31 && x == 22) || (y == 32 && x == 22) || (y == 33 && x == 22) || (y == 47 && x == 22) || (y == 48 && x == 22) || (y == 49 && x == 22) || (y == 50 && x == 22) || (y == 51 && x == 22) || (y == 52 && x == 22) || (y == 53 && x == 22) || (y == 54 && x == 22) || (y == 55 && x == 22) || (y == 56 && x == 22) || (y == 57 && x == 22) || (y == 58 && x == 22) || (y == 59 && x == 22) || (y == 60 && x == 22) || (y == 61 && x == 22) || (y == 62 && x == 22) || (y == 63 && x == 22) || (y == 0 && x == 23) || (y == 1 && x == 23) || (y == 2 && x == 23) || (y == 3 && x == 23) || (y == 4 && x == 23) || (y == 5 && x == 23) || (y == 6 && x == 23) || (y == 7 && x == 23) || (y == 8 && x == 23) || (y == 9 && x == 23) || (y == 10 && x == 23) || (y == 11 && x == 23) || (y == 12 && x == 23) || (y == 13 && x == 23) || (y == 14 && x == 23) || (y == 15 && x == 23) || (y == 16 && x == 23) || (y == 17 && x == 23) || (y == 18 && x == 23) || (y == 19 && x == 23) || (y == 20 && x == 23) || (y == 21 && x == 23) || (y == 22 && x == 23) || (y == 23 && x == 23) || (y == 24 && x == 23) || (y == 25 && x == 23) || (y == 26 && x == 23) || (y == 27 && x == 23) || (y == 28 && x == 23) || (y == 29 && x == 23) || (y == 30 && x == 23) || (y == 31 && x == 23) || (y == 49 && x == 23) || (y == 50 && x == 23) || (y == 51 && x == 23) || (y == 52 && x == 23) || (y == 53 && x == 23) || (y == 54 && x == 23) || (y == 55 && x == 23) || (y == 56 && x == 23) || (y == 57 && x == 23) || (y == 58 && x == 23) || (y == 59 && x == 23) || (y == 60 && x == 23) || (y == 61 && x == 23) || (y == 62 && x == 23) || (y == 63 && x == 23) || (y == 0 && x == 24) || (y == 1 && x == 24) || (y == 2 && x == 24) || (y == 3 && x == 24) || (y == 4 && x == 24) || (y == 5 && x == 24) || (y == 6 && x == 24) || (y == 7 && x == 24) || (y == 8 && x == 24) || (y == 9 && x == 24) || (y == 10 && x == 24) || (y == 11 && x == 24) || (y == 12 && x == 24) || (y == 13 && x == 24) || (y == 14 && x == 24) || (y == 15 && x == 24) || (y == 16 && x == 24) || (y == 17 && x == 24) || (y == 18 && x == 24) || (y == 19 && x == 24) || (y == 20 && x == 24) || (y == 21 && x == 24) || (y == 22 && x == 24) || (y == 23 && x == 24) || (y == 24 && x == 24) || (y == 25 && x == 24) || (y == 26 && x == 24) || (y == 27 && x == 24) || (y == 28 && x == 24) || (y == 29 && x == 24) || (y == 30 && x == 24) || (y == 50 && x == 24) || (y == 51 && x == 24) || (y == 52 && x == 24) || (y == 53 && x == 24) || (y == 54 && x == 24) || (y == 55 && x == 24) || (y == 56 && x == 24) || (y == 57 && x == 24) || (y == 58 && x == 24) || (y == 59 && x == 24) || (y == 60 && x == 24) || (y == 61 && x == 24) || (y == 62 && x == 24) || (y == 63 && x == 24) || (y == 0 && x == 25) || (y == 1 && x == 25) || (y == 2 && x == 25) || (y == 3 && x == 25) || (y == 4 && x == 25) || (y == 5 && x == 25) || (y == 6 && x == 25) || (y == 7 && x == 25) || (y == 8 && x == 25) || (y == 9 && x == 25) || (y == 10 && x == 25) || (y == 11 && x == 25) || (y == 12 && x == 25) || (y == 13 && x == 25) || (y == 14 && x == 25) || (y == 15 && x == 25) || (y == 16 && x == 25) || (y == 17 && x == 25) || (y == 18 && x == 25) || (y == 19 && x == 25) || (y == 20 && x == 25) || (y == 21 && x == 25) || (y == 22 && x == 25) || (y == 23 && x == 25) || (y == 24 && x == 25) || (y == 25 && x == 25) || (y == 26 && x == 25) || (y == 27 && x == 25) || (y == 28 && x == 25) || (y == 29 && x == 25) || (y == 51 && x == 25) || (y == 52 && x == 25) || (y == 53 && x == 25) || (y == 54 && x == 25) || (y == 55 && x == 25) || (y == 56 && x == 25) || (y == 57 && x == 25) || (y == 58 && x == 25) || (y == 59 && x == 25) || (y == 60 && x == 25) || (y == 61 && x == 25) || (y == 62 && x == 25) || (y == 63 && x == 25) || (y == 0 && x == 26) || (y == 1 && x == 26) || (y == 2 && x == 26) || (y == 3 && x == 26) || (y == 4 && x == 26) || (y == 5 && x == 26) || (y == 6 && x == 26) || (y == 7 && x == 26) || (y == 8 && x == 26) || (y == 9 && x == 26) || (y == 10 && x == 26) || (y == 11 && x == 26) || (y == 12 && x == 26) || (y == 13 && x == 26) || (y == 14 && x == 26) || (y == 15 && x == 26) || (y == 16 && x == 26) || (y == 17 && x == 26) || (y == 18 && x == 26) || (y == 19 && x == 26) || (y == 20 && x == 26) || (y == 21 && x == 26) || (y == 22 && x == 26) || (y == 23 && x == 26) || (y == 24 && x == 26) || (y == 25 && x == 26) || (y == 26 && x == 26) || (y == 27 && x == 26) || (y == 28 && x == 26) || (y == 53 && x == 26) || (y == 54 && x == 26) || (y == 55 && x == 26) || (y == 56 && x == 26) || (y == 57 && x == 26) || (y == 58 && x == 26) || (y == 59 && x == 26) || (y == 60 && x == 26) || (y == 61 && x == 26) || (y == 62 && x == 26) || (y == 63 && x == 26) || (y == 0 && x == 27) || (y == 1 && x == 27) || (y == 2 && x == 27) || (y == 3 && x == 27) || (y == 4 && x == 27) || (y == 5 && x == 27) || (y == 6 && x == 27) || (y == 7 && x == 27) || (y == 8 && x == 27) || (y == 9 && x == 27) || (y == 10 && x == 27) || (y == 11 && x == 27) || (y == 12 && x == 27) || (y == 13 && x == 27) || (y == 14 && x == 27) || (y == 15 && x == 27) || (y == 16 && x == 27) || (y == 17 && x == 27) || (y == 18 && x == 27) || (y == 19 && x == 27) || (y == 20 && x == 27) || (y == 21 && x == 27) || (y == 22 && x == 27) || (y == 23 && x == 27) || (y == 24 && x == 27) || (y == 25 && x == 27) || (y == 26 && x == 27) || (y == 54 && x == 27) || (y == 55 && x == 27) || (y == 56 && x == 27) || (y == 57 && x == 27) || (y == 58 && x == 27) || (y == 59 && x == 27) || (y == 60 && x == 27) || (y == 61 && x == 27) || (y == 62 && x == 27) || (y == 63 && x == 27) || (y == 0 && x == 28) || (y == 1 && x == 28) || (y == 2 && x == 28) || (y == 3 && x == 28) || (y == 4 && x == 28) || (y == 5 && x == 28) || (y == 6 && x == 28) || (y == 7 && x == 28) || (y == 8 && x == 28) || (y == 9 && x == 28) || (y == 10 && x == 28) || (y == 11 && x == 28) || (y == 12 && x == 28) || (y == 13 && x == 28) || (y == 14 && x == 28) || (y == 15 && x == 28) || (y == 16 && x == 28) || (y == 17 && x == 28) || (y == 18 && x == 28) || (y == 19 && x == 28) || (y == 20 && x == 28) || (y == 21 && x == 28) || (y == 22 && x == 28) || (y == 23 && x == 28) || (y == 24 && x == 28) || (y == 25 && x == 28) || (y == 26 && x == 28) || (y == 55 && x == 28) || (y == 56 && x == 28) || (y == 57 && x == 28) || (y == 58 && x == 28) || (y == 59 && x == 28) || (y == 60 && x == 28) || (y == 61 && x == 28) || (y == 62 && x == 28) || (y == 63 && x == 28) || (y == 0 && x == 29) || (y == 1 && x == 29) || (y == 2 && x == 29) || (y == 3 && x == 29) || (y == 4 && x == 29) || (y == 5 && x == 29) || (y == 6 && x == 29) || (y == 7 && x == 29) || (y == 8 && x == 29) || (y == 9 && x == 29) || (y == 10 && x == 29) || (y == 11 && x == 29) || (y == 12 && x == 29) || (y == 13 && x == 29) || (y == 14 && x == 29) || (y == 15 && x == 29) || (y == 16 && x == 29) || (y == 17 && x == 29) || (y == 18 && x == 29) || (y == 19 && x == 29) || (y == 20 && x == 29) || (y == 21 && x == 29) || (y == 22 && x == 29) || (y == 23 && x == 29) || (y == 24 && x == 29) || (y == 55 && x == 29) || (y == 56 && x == 29) || (y == 57 && x == 29) || (y == 58 && x == 29) || (y == 59 && x == 29) || (y == 60 && x == 29) || (y == 61 && x == 29) || (y == 62 && x == 29) || (y == 63 && x == 29) || (y == 0 && x == 30) || (y == 1 && x == 30) || (y == 2 && x == 30) || (y == 3 && x == 30) || (y == 4 && x == 30) || (y == 5 && x == 30) || (y == 6 && x == 30) || (y == 7 && x == 30) || (y == 8 && x == 30) || (y == 9 && x == 30) || (y == 10 && x == 30) || (y == 11 && x == 30) || (y == 12 && x == 30) || (y == 13 && x == 30) || (y == 14 && x == 30) || (y == 15 && x == 30) || (y == 16 && x == 30) || (y == 17 && x == 30) || (y == 18 && x == 30) || (y == 19 && x == 30) || (y == 20 && x == 30) || (y == 21 && x == 30) || (y == 22 && x == 30) || (y == 56 && x == 30) || (y == 57 && x == 30) || (y == 58 && x == 30) || (y == 59 && x == 30) || (y == 60 && x == 30) || (y == 61 && x == 30) || (y == 62 && x == 30) || (y == 63 && x == 30) || (y == 0 && x == 31) || (y == 1 && x == 31) || (y == 2 && x == 31) || (y == 13 && x == 31) || (y == 14 && x == 31) || (y == 15 && x == 31) || (y == 16 && x == 31) || (y == 17 && x == 31) || (y == 18 && x == 31) || (y == 19 && x == 31) || (y == 20 && x == 31) || (y == 21 && x == 31) || (y == 57 && x == 31) || (y == 58 && x == 31) || (y == 59 && x == 31) || (y == 60 && x == 31) || (y == 61 && x == 31) || (y == 62 && x == 31) || (y == 63 && x == 31) || (y == 0 && x == 32) || (y == 1 && x == 32) || (y == 2 && x == 32) || (y == 13 && x == 32) || (y == 14 && x == 32) || (y == 15 && x == 32) || (y == 16 && x == 32) || (y == 17 && x == 32) || (y == 18 && x == 32) || (y == 19 && x == 32) || (y == 57 && x == 32) || (y == 58 && x == 32) || (y == 59 && x == 32) || (y == 60 && x == 32) || (y == 61 && x == 32) || (y == 62 && x == 32) || (y == 63 && x == 32) || (y == 0 && x == 33) || (y == 1 && x == 33) || (y == 2 && x == 33) || (y == 3 && x == 33) || (y == 4 && x == 33) || (y == 5 && x == 33) || (y == 6 && x == 33) || (y == 7 && x == 33) || (y == 8 && x == 33) || (y == 9 && x == 33) || (y == 10 && x == 33) || (y == 13 && x == 33) || (y == 14 && x == 33) || (y == 15 && x == 33) || (y == 16 && x == 33) || (y == 17 && x == 33) || (y == 18 && x == 33) || (y == 58 && x == 33) || (y == 59 && x == 33) || (y == 60 && x == 33) || (y == 61 && x == 33) || (y == 62 && x == 33) || (y == 63 && x == 33) || (y == 0 && x == 34) || (y == 1 && x == 34) || (y == 2 && x == 34) || (y == 3 && x == 34) || (y == 4 && x == 34) || (y == 5 && x == 34) || (y == 6 && x == 34) || (y == 7 && x == 34) || (y == 8 && x == 34) || (y == 9 && x == 34) || (y == 10 && x == 34) || (y == 13 && x == 34) || (y == 14 && x == 34) || (y == 15 && x == 34) || (y == 16 && x == 34) || (y == 17 && x == 34) || (y == 58 && x == 34) || (y == 59 && x == 34) || (y == 60 && x == 34) || (y == 61 && x == 34) || (y == 62 && x == 34) || (y == 63 && x == 34) || (y == 0 && x == 35) || (y == 1 && x == 35) || (y == 2 && x == 35) || (y == 3 && x == 35) || (y == 4 && x == 35) || (y == 5 && x == 35) || (y == 6 && x == 35) || (y == 7 && x == 35) || (y == 8 && x == 35) || (y == 9 && x == 35) || (y == 10 && x == 35) || (y == 13 && x == 35) || (y == 14 && x == 35) || (y == 15 && x == 35) || (y == 16 && x == 35) || (y == 17 && x == 35) || (y == 58 && x == 35) || (y == 59 && x == 35) || (y == 60 && x == 35) || (y == 61 && x == 35) || (y == 62 && x == 35) || (y == 63 && x == 35) || (y == 0 && x == 36) || (y == 1 && x == 36) || (y == 2 && x == 36) || (y == 3 && x == 36) || (y == 4 && x == 36) || (y == 5 && x == 36) || (y == 6 && x == 36) || (y == 7 && x == 36) || (y == 8 && x == 36) || (y == 9 && x == 36) || (y == 10 && x == 36) || (y == 13 && x == 36) || (y == 14 && x == 36) || (y == 15 && x == 36) || (y == 16 && x == 36) || (y == 58 && x == 36) || (y == 59 && x == 36) || (y == 60 && x == 36) || (y == 61 && x == 36) || (y == 62 && x == 36) || (y == 63 && x == 36) || (y == 0 && x == 37) || (y == 1 && x == 37) || (y == 2 && x == 37) || (y == 3 && x == 37) || (y == 4 && x == 37) || (y == 5 && x == 37) || (y == 6 && x == 37) || (y == 7 && x == 37) || (y == 8 && x == 37) || (y == 9 && x == 37) || (y == 10 && x == 37) || (y == 13 && x == 37) || (y == 14 && x == 37) || (y == 15 && x == 37) || (y == 16 && x == 37) || (y == 58 && x == 37) || (y == 59 && x == 37) || (y == 60 && x == 37) || (y == 61 && x == 37) || (y == 62 && x == 37) || (y == 63 && x == 37) || (y == 0 && x == 38) || (y == 1 && x == 38) || (y == 2 && x == 38) || (y == 3 && x == 38) || (y == 4 && x == 38) || (y == 5 && x == 38) || (y == 6 && x == 38) || (y == 7 && x == 38) || (y == 8 && x == 38) || (y == 9 && x == 38) || (y == 10 && x == 38) || (y == 13 && x == 38) || (y == 14 && x == 38) || (y == 15 && x == 38) || (y == 58 && x == 38) || (y == 59 && x == 38) || (y == 60 && x == 38) || (y == 61 && x == 38) || (y == 62 && x == 38) || (y == 63 && x == 38) || (y == 0 && x == 39) || (y == 1 && x == 39) || (y == 2 && x == 39) || (y == 3 && x == 39) || (y == 4 && x == 39) || (y == 5 && x == 39) || (y == 6 && x == 39) || (y == 7 && x == 39) || (y == 8 && x == 39) || (y == 9 && x == 39) || (y == 10 && x == 39) || (y == 11 && x == 39) || (y == 12 && x == 39) || (y == 13 && x == 39) || (y == 14 && x == 39) || (y == 15 && x == 39) || (y == 58 && x == 39) || (y == 59 && x == 39) || (y == 60 && x == 39) || (y == 61 && x == 39) || (y == 62 && x == 39) || (y == 63 && x == 39) || (y == 0 && x == 40) || (y == 1 && x == 40) || (y == 2 && x == 40) || (y == 3 && x == 40) || (y == 4 && x == 40) || (y == 5 && x == 40) || (y == 6 && x == 40) || (y == 7 && x == 40) || (y == 8 && x == 40) || (y == 9 && x == 40) || (y == 10 && x == 40) || (y == 11 && x == 40) || (y == 12 && x == 40) || (y == 13 && x == 40) || (y == 14 && x == 40) || (y == 15 && x == 40) || (y == 58 && x == 40) || (y == 0 && x == 41) || (y == 1 && x == 41) || (y == 2 && x == 41) || (y == 13 && x == 41) || (y == 14 && x == 41) || (y == 15 && x == 41) || (y == 57 && x == 41) || (y == 58 && x == 41) || (y == 60 && x == 41) || (y == 63 && x == 41) || (y == 0 && x == 42) || (y == 1 && x == 42) || (y == 2 && x == 42) || (y == 13 && x == 42) || (y == 14 && x == 42) || (y == 15 && x == 42) || (y == 57 && x == 42) || (y == 58 && x == 42) || (y == 62 && x == 42) || (y == 0 && x == 43) || (y == 1 && x == 43) || (y == 2 && x == 43) || (y == 5 && x == 43) || (y == 6 && x == 43) || (y == 7 && x == 43) || (y == 8 && x == 43) || (y == 9 && x == 43) || (y == 10 && x == 43) || (y == 13 && x == 43) || (y == 14 && x == 43) || (y == 15 && x == 43) || (y == 57 && x == 43) || (y == 58 && x == 43) || (y == 59 && x == 43) || (y == 60 && x == 43) || (y == 61 && x == 43) || (y == 62 && x == 43) || (y == 63 && x == 43) || (y == 0 && x == 44) || (y == 1 && x == 44) || (y == 2 && x == 44) || (y == 5 && x == 44) || (y == 6 && x == 44) || (y == 7 && x == 44) || (y == 8 && x == 44) || (y == 9 && x == 44) || (y == 10 && x == 44) || (y == 13 && x == 44) || (y == 14 && x == 44) || (y == 15 && x == 44) || (y == 57 && x == 44) || (y == 58 && x == 44) || (y == 0 && x == 45) || (y == 1 && x == 45) || (y == 2 && x == 45) || (y == 5 && x == 45) || (y == 6 && x == 45) || (y == 7 && x == 45) || (y == 8 && x == 45) || (y == 9 && x == 45) || (y == 10 && x == 45) || (y == 13 && x == 45) || (y == 14 && x == 45) || (y == 57 && x == 45) || (y == 58 && x == 45) || (y == 60 && x == 45) || (y == 62 && x == 45) || (y == 0 && x == 46) || (y == 1 && x == 46) || (y == 2 && x == 46) || (y == 5 && x == 46) || (y == 6 && x == 46) || (y == 7 && x == 46) || (y == 8 && x == 46) || (y == 9 && x == 46) || (y == 10 && x == 46) || (y == 13 && x == 46) || (y == 14 && x == 46) || (y == 57 && x == 46) || (y == 58 && x == 46) || (y == 60 && x == 46) || (y == 62 && x == 46) || (y == 0 && x == 47) || (y == 1 && x == 47) || (y == 2 && x == 47) || (y == 13 && x == 47) || (y == 14 && x == 47) || (y == 58 && x == 47) || (y == 59 && x == 47) || (y == 60 && x == 47) || (y == 61 && x == 47) || (y == 62 && x == 47) || (y == 63 && x == 47) || (y == 0 && x == 48) || (y == 1 && x == 48) || (y == 2 && x == 48) || (y == 13 && x == 48) || (y == 14 && x == 48) || (y == 58 && x == 48) || (y == 62 && x == 48) || (y == 0 && x == 49) || (y == 1 && x == 49) || (y == 2 && x == 49) || (y == 3 && x == 49) || (y == 4 && x == 49) || (y == 5 && x == 49) || (y == 6 && x == 49) || (y == 7 && x == 49) || (y == 8 && x == 49) || (y == 9 && x == 49) || (y == 10 && x == 49) || (y == 11 && x == 49) || (y == 12 && x == 49) || (y == 13 && x == 49) || (y == 14 && x == 49) || (y == 58 && x == 49) || (y == 60 && x == 49) || (y == 62 && x == 49) || (y == 0 && x == 50) || (y == 1 && x == 50) || (y == 2 && x == 50) || (y == 3 && x == 50) || (y == 4 && x == 50) || (y == 5 && x == 50) || (y == 6 && x == 50) || (y == 7 && x == 50) || (y == 8 && x == 50) || (y == 9 && x == 50) || (y == 10 && x == 50) || (y == 11 && x == 50) || (y == 12 && x == 50) || (y == 13 && x == 50) || (y == 14 && x == 50) || (y == 58 && x == 50) || (y == 60 && x == 50) || (y == 0 && x == 51) || (y == 1 && x == 51) || (y == 2 && x == 51) || (y == 13 && x == 51) || (y == 14 && x == 51) || (y == 58 && x == 51) || (y == 59 && x == 51) || (y == 60 && x == 51) || (y == 61 && x == 51) || (y == 62 && x == 51) || (y == 63 && x == 51) || (y == 0 && x == 52) || (y == 1 && x == 52) || (y == 2 && x == 52) || (y == 13 && x == 52) || (y == 14 && x == 52) || (y == 57 && x == 52) || (y == 58 && x == 52) || (y == 0 && x == 53) || (y == 1 && x == 53) || (y == 2 && x == 53) || (y == 5 && x == 53) || (y == 6 && x == 53) || (y == 9 && x == 53) || (y == 10 && x == 53) || (y == 13 && x == 53) || (y == 14 && x == 53) || (y == 57 && x == 53) || (y == 58 && x == 53) || (y == 60 && x == 53) || (y == 62 && x == 53) || (y == 0 && x == 54) || (y == 1 && x == 54) || (y == 2 && x == 54) || (y == 5 && x == 54) || (y == 6 && x == 54) || (y == 9 && x == 54) || (y == 10 && x == 54) || (y == 13 && x == 54) || (y == 14 && x == 54) || (y == 57 && x == 54) || (y == 58 && x == 54) || (y == 60 && x == 54) || (y == 62 && x == 54) || (y == 0 && x == 55) || (y == 1 && x == 55) || (y == 2 && x == 55) || (y == 5 && x == 55) || (y == 6 && x == 55) || (y == 9 && x == 55) || (y == 10 && x == 55) || (y == 13 && x == 55) || (y == 14 && x == 55) || (y == 57 && x == 55) || (y == 58 && x == 55) || (y == 59 && x == 55) || (y == 60 && x == 55) || (y == 61 && x == 55) || (y == 62 && x == 55) || (y == 63 && x == 55) || (y == 0 && x == 56) || (y == 1 && x == 56) || (y == 2 && x == 56) || (y == 5 && x == 56) || (y == 6 && x == 56) || (y == 9 && x == 56) || (y == 10 && x == 56) || (y == 13 && x == 56) || (y == 14 && x == 56) || (y == 57 && x == 56) || (y == 58 && x == 56) || (y == 60 && x == 56) || (y == 61 && x == 56) || (y == 62 && x == 56) || (y == 63 && x == 56) || (y == 0 && x == 57) || (y == 1 && x == 57) || (y == 2 && x == 57) || (y == 5 && x == 57) || (y == 6 && x == 57) || (y == 13 && x == 57) || (y == 14 && x == 57) || (y == 15 && x == 57) || (y == 57 && x == 57) || (y == 58 && x == 57) || (y == 0 && x == 58) || (y == 1 && x == 58) || (y == 2 && x == 58) || (y == 5 && x == 58) || (y == 6 && x == 58) || (y == 13 && x == 58) || (y == 14 && x == 58) || (y == 15 && x == 58) || (y == 57 && x == 58) || (y == 58 && x == 58) || (y == 60 && x == 58) || (y == 61 && x == 58) || (y == 62 && x == 58) || (y == 63 && x == 58) || (y == 0 && x == 59) || (y == 1 && x == 59) || (y == 2 && x == 59) || (y == 3 && x == 59) || (y == 4 && x == 59) || (y == 5 && x == 59) || (y == 6 && x == 59) || (y == 7 && x == 59) || (y == 8 && x == 59) || (y == 9 && x == 59) || (y == 10 && x == 59) || (y == 11 && x == 59) || (y == 12 && x == 59) || (y == 13 && x == 59) || (y == 14 && x == 59) || (y == 15 && x == 59) || (y == 56 && x == 59) || (y == 57 && x == 59) || (y == 58 && x == 59) || (y == 59 && x == 59) || (y == 60 && x == 59) || (y == 61 && x == 59) || (y == 62 && x == 59) || (y == 63 && x == 59) || (y == 0 && x == 60) || (y == 1 && x == 60) || (y == 2 && x == 60) || (y == 3 && x == 60) || (y == 4 && x == 60) || (y == 5 && x == 60) || (y == 6 && x == 60) || (y == 7 && x == 60) || (y == 8 && x == 60) || (y == 9 && x == 60) || (y == 10 && x == 60) || (y == 11 && x == 60) || (y == 12 && x == 60) || (y == 13 && x == 60) || (y == 14 && x == 60) || (y == 15 && x == 60) || (y == 16 && x == 60) || (y == 56 && x == 60) || (y == 57 && x == 60) || (y == 58 && x == 60) || (y == 59 && x == 60) || (y == 60 && x == 60) || (y == 61 && x == 60) || (y == 62 && x == 60) || (y == 63 && x == 60) || (y == 0 && x == 61) || (y == 1 && x == 61) || (y == 2 && x == 61) || (y == 13 && x == 61) || (y == 14 && x == 61) || (y == 15 && x == 61) || (y == 16 && x == 61) || (y == 17 && x == 61) || (y == 56 && x == 61) || (y == 57 && x == 61) || (y == 58 && x == 61) || (y == 59 && x == 61) || (y == 60 && x == 61) || (y == 61 && x == 61) || (y == 62 && x == 61) || (y == 63 && x == 61) || (y == 0 && x == 62) || (y == 1 && x == 62) || (y == 2 && x == 62) || (y == 13 && x == 62) || (y == 14 && x == 62) || (y == 15 && x == 62) || (y == 16 && x == 62) || (y == 17 && x == 62) || (y == 18 && x == 62) || (y == 55 && x == 62) || (y == 56 && x == 62) || (y == 57 && x == 62) || (y == 58 && x == 62) || (y == 59 && x == 62) || (y == 60 && x == 62) || (y == 61 && x == 62) || (y == 62 && x == 62) || (y == 63 && x == 62) || (y == 0 && x == 63) || (y == 1 && x == 63) || (y == 2 && x == 63) || (y == 5 && x == 63) || (y == 6 && x == 63) || (y == 9 && x == 63) || (y == 10 && x == 63) || (y == 13 && x == 63) || (y == 14 && x == 63) || (y == 15 && x == 63) || (y == 16 && x == 63) || (y == 17 && x == 63) || (y == 18 && x == 63) || (y == 19 && x == 63) || (y == 55 && x == 63) || (y == 56 && x == 63) || (y == 57 && x == 63) || (y == 58 && x == 63) || (y == 59 && x == 63) || (y == 60 && x == 63) || (y == 61 && x == 63) || (y == 62 && x == 63) || (y == 63 && x == 63) || (y == 0 && x == 64) || (y == 1 && x == 64) || (y == 2 && x == 64) || (y == 5 && x == 64) || (y == 6 && x == 64) || (y == 9 && x == 64) || (y == 10 && x == 64) || (y == 13 && x == 64) || (y == 14 && x == 64) || (y == 15 && x == 64) || (y == 16 && x == 64) || (y == 17 && x == 64) || (y == 18 && x == 64) || (y == 19 && x == 64) || (y == 20 && x == 64) || (y == 55 && x == 64) || (y == 56 && x == 64) || (y == 57 && x == 64) || (y == 58 && x == 64) || (y == 59 && x == 64) || (y == 60 && x == 64) || (y == 61 && x == 64) || (y == 62 && x == 64) || (y == 63 && x == 64) || (y == 0 && x == 65) || (y == 1 && x == 65) || (y == 2 && x == 65) || (y == 5 && x == 65) || (y == 6 && x == 65) || (y == 9 && x == 65) || (y == 10 && x == 65) || (y == 13 && x == 65) || (y == 14 && x == 65) || (y == 15 && x == 65) || (y == 16 && x == 65) || (y == 17 && x == 65) || (y == 18 && x == 65) || (y == 19 && x == 65) || (y == 20 && x == 65) || (y == 21 && x == 65) || (y == 54 && x == 65) || (y == 55 && x == 65) || (y == 56 && x == 65) || (y == 57 && x == 65) || (y == 58 && x == 65) || (y == 59 && x == 65) || (y == 60 && x == 65) || (y == 61 && x == 65) || (y == 62 && x == 65) || (y == 63 && x == 65) || (y == 0 && x == 66) || (y == 1 && x == 66) || (y == 2 && x == 66) || (y == 5 && x == 66) || (y == 6 && x == 66) || (y == 9 && x == 66) || (y == 10 && x == 66) || (y == 13 && x == 66) || (y == 14 && x == 66) || (y == 15 && x == 66) || (y == 16 && x == 66) || (y == 17 && x == 66) || (y == 18 && x == 66) || (y == 19 && x == 66) || (y == 20 && x == 66) || (y == 21 && x == 66) || (y == 22 && x == 66) || (y == 54 && x == 66) || (y == 55 && x == 66) || (y == 56 && x == 66) || (y == 57 && x == 66) || (y == 58 && x == 66) || (y == 59 && x == 66) || (y == 60 && x == 66) || (y == 61 && x == 66) || (y == 62 && x == 66) || (y == 63 && x == 66) || (y == 0 && x == 67) || (y == 1 && x == 67) || (y == 2 && x == 67) || (y == 5 && x == 67) || (y == 6 && x == 67) || (y == 9 && x == 67) || (y == 10 && x == 67) || (y == 13 && x == 67) || (y == 14 && x == 67) || (y == 15 && x == 67) || (y == 16 && x == 67) || (y == 17 && x == 67) || (y == 18 && x == 67) || (y == 19 && x == 67) || (y == 20 && x == 67) || (y == 21 && x == 67) || (y == 22 && x == 67) || (y == 23 && x == 67) || (y == 54 && x == 67) || (y == 55 && x == 67) || (y == 56 && x == 67) || (y == 57 && x == 67) || (y == 58 && x == 67) || (y == 59 && x == 67) || (y == 60 && x == 67) || (y == 61 && x == 67) || (y == 62 && x == 67) || (y == 63 && x == 67) || (y == 0 && x == 68) || (y == 1 && x == 68) || (y == 2 && x == 68) || (y == 5 && x == 68) || (y == 6 && x == 68) || (y == 9 && x == 68) || (y == 10 && x == 68) || (y == 13 && x == 68) || (y == 14 && x == 68) || (y == 15 && x == 68) || (y == 16 && x == 68) || (y == 17 && x == 68) || (y == 18 && x == 68) || (y == 19 && x == 68) || (y == 20 && x == 68) || (y == 21 && x == 68) || (y == 22 && x == 68) || (y == 23 && x == 68) || (y == 24 && x == 68) || (y == 53 && x == 68) || (y == 54 && x == 68) || (y == 55 && x == 68) || (y == 56 && x == 68) || (y == 57 && x == 68) || (y == 58 && x == 68) || (y == 59 && x == 68) || (y == 60 && x == 68) || (y == 61 && x == 68) || (y == 62 && x == 68) || (y == 63 && x == 68) || (y == 0 && x == 69) || (y == 1 && x == 69) || (y == 2 && x == 69) || (y == 3 && x == 69) || (y == 4 && x == 69) || (y == 5 && x == 69) || (y == 6 && x == 69) || (y == 7 && x == 69) || (y == 8 && x == 69) || (y == 9 && x == 69) || (y == 10 && x == 69) || (y == 11 && x == 69) || (y == 12 && x == 69) || (y == 13 && x == 69) || (y == 14 && x == 69) || (y == 15 && x == 69) || (y == 16 && x == 69) || (y == 17 && x == 69) || (y == 18 && x == 69) || (y == 19 && x == 69) || (y == 20 && x == 69) || (y == 21 && x == 69) || (y == 22 && x == 69) || (y == 23 && x == 69) || (y == 24 && x == 69) || (y == 25 && x == 69) || (y == 53 && x == 69) || (y == 54 && x == 69) || (y == 55 && x == 69) || (y == 56 && x == 69) || (y == 57 && x == 69) || (y == 58 && x == 69) || (y == 59 && x == 69) || (y == 60 && x == 69) || (y == 61 && x == 69) || (y == 62 && x == 69) || (y == 63 && x == 69) || (y == 0 && x == 70) || (y == 1 && x == 70) || (y == 2 && x == 70) || (y == 3 && x == 70) || (y == 4 && x == 70) || (y == 5 && x == 70) || (y == 6 && x == 70) || (y == 7 && x == 70) || (y == 8 && x == 70) || (y == 9 && x == 70) || (y == 10 && x == 70) || (y == 11 && x == 70) || (y == 12 && x == 70) || (y == 13 && x == 70) || (y == 14 && x == 70) || (y == 15 && x == 70) || (y == 16 && x == 70) || (y == 17 && x == 70) || (y == 18 && x == 70) || (y == 19 && x == 70) || (y == 20 && x == 70) || (y == 21 && x == 70) || (y == 22 && x == 70) || (y == 23 && x == 70) || (y == 24 && x == 70) || (y == 25 && x == 70) || (y == 26 && x == 70) || (y == 52 && x == 70) || (y == 53 && x == 70) || (y == 54 && x == 70) || (y == 55 && x == 70) || (y == 56 && x == 70) || (y == 57 && x == 70) || (y == 58 && x == 70) || (y == 59 && x == 70) || (y == 60 && x == 70) || (y == 61 && x == 70) || (y == 62 && x == 70) || (y == 63 && x == 70) || (y == 0 && x == 71) || (y == 1 && x == 71) || (y == 2 && x == 71) || (y == 3 && x == 71) || (y == 4 && x == 71) || (y == 5 && x == 71) || (y == 6 && x == 71) || (y == 7 && x == 71) || (y == 8 && x == 71) || (y == 9 && x == 71) || (y == 10 && x == 71) || (y == 11 && x == 71) || (y == 12 && x == 71) || (y == 13 && x == 71) || (y == 14 && x == 71) || (y == 15 && x == 71) || (y == 16 && x == 71) || (y == 17 && x == 71) || (y == 18 && x == 71) || (y == 19 && x == 71) || (y == 20 && x == 71) || (y == 21 && x == 71) || (y == 22 && x == 71) || (y == 23 && x == 71) || (y == 24 && x == 71) || (y == 25 && x == 71) || (y == 26 && x == 71) || (y == 27 && x == 71) || (y == 28 && x == 71) || (y == 51 && x == 71) || (y == 52 && x == 71) || (y == 53 && x == 71) || (y == 54 && x == 71) || (y == 55 && x == 71) || (y == 56 && x == 71) || (y == 57 && x == 71) || (y == 58 && x == 71) || (y == 59 && x == 71) || (y == 60 && x == 71) || (y == 61 && x == 71) || (y == 62 && x == 71) || (y == 63 && x == 71) || (y == 0 && x == 72) || (y == 1 && x == 72) || (y == 2 && x == 72) || (y == 3 && x == 72) || (y == 4 && x == 72) || (y == 5 && x == 72) || (y == 6 && x == 72) || (y == 7 && x == 72) || (y == 8 && x == 72) || (y == 9 && x == 72) || (y == 10 && x == 72) || (y == 11 && x == 72) || (y == 12 && x == 72) || (y == 13 && x == 72) || (y == 14 && x == 72) || (y == 15 && x == 72) || (y == 16 && x == 72) || (y == 17 && x == 72) || (y == 18 && x == 72) || (y == 19 && x == 72) || (y == 20 && x == 72) || (y == 21 && x == 72) || (y == 22 && x == 72) || (y == 23 && x == 72) || (y == 24 && x == 72) || (y == 25 && x == 72) || (y == 26 && x == 72) || (y == 27 && x == 72) || (y == 28 && x == 72) || (y == 29 && x == 72) || (y == 50 && x == 72) || (y == 51 && x == 72) || (y == 52 && x == 72) || (y == 53 && x == 72) || (y == 54 && x == 72) || (y == 55 && x == 72) || (y == 56 && x == 72) || (y == 57 && x == 72) || (y == 58 && x == 72) || (y == 59 && x == 72) || (y == 60 && x == 72) || (y == 61 && x == 72) || (y == 62 && x == 72) || (y == 63 && x == 72) || (y == 0 && x == 73) || (y == 1 && x == 73) || (y == 2 && x == 73) || (y == 3 && x == 73) || (y == 4 && x == 73) || (y == 5 && x == 73) || (y == 6 && x == 73) || (y == 7 && x == 73) || (y == 8 && x == 73) || (y == 9 && x == 73) || (y == 10 && x == 73) || (y == 11 && x == 73) || (y == 12 && x == 73) || (y == 13 && x == 73) || (y == 14 && x == 73) || (y == 15 && x == 73) || (y == 16 && x == 73) || (y == 17 && x == 73) || (y == 18 && x == 73) || (y == 19 && x == 73) || (y == 20 && x == 73) || (y == 21 && x == 73) || (y == 22 && x == 73) || (y == 23 && x == 73) || (y == 24 && x == 73) || (y == 25 && x == 73) || (y == 26 && x == 73) || (y == 27 && x == 73) || (y == 28 && x == 73) || (y == 29 && x == 73) || (y == 30 && x == 73) || (y == 49 && x == 73) || (y == 50 && x == 73) || (y == 51 && x == 73) || (y == 52 && x == 73) || (y == 53 && x == 73) || (y == 54 && x == 73) || (y == 55 && x == 73) || (y == 56 && x == 73) || (y == 57 && x == 73) || (y == 58 && x == 73) || (y == 59 && x == 73) || (y == 60 && x == 73) || (y == 61 && x == 73) || (y == 62 && x == 73) || (y == 63 && x == 73) || (y == 0 && x == 74) || (y == 1 && x == 74) || (y == 2 && x == 74) || (y == 3 && x == 74) || (y == 4 && x == 74) || (y == 5 && x == 74) || (y == 6 && x == 74) || (y == 7 && x == 74) || (y == 8 && x == 74) || (y == 9 && x == 74) || (y == 10 && x == 74) || (y == 11 && x == 74) || (y == 12 && x == 74) || (y == 13 && x == 74) || (y == 14 && x == 74) || (y == 15 && x == 74) || (y == 16 && x == 74) || (y == 17 && x == 74) || (y == 18 && x == 74) || (y == 19 && x == 74) || (y == 20 && x == 74) || (y == 21 && x == 74) || (y == 22 && x == 74) || (y == 23 && x == 74) || (y == 24 && x == 74) || (y == 25 && x == 74) || (y == 26 && x == 74) || (y == 27 && x == 74) || (y == 28 && x == 74) || (y == 29 && x == 74) || (y == 30 && x == 74) || (y == 31 && x == 74) || (y == 32 && x == 74) || (y == 47 && x == 74) || (y == 48 && x == 74) || (y == 49 && x == 74) || (y == 50 && x == 74) || (y == 51 && x == 74) || (y == 52 && x == 74) || (y == 53 && x == 74) || (y == 54 && x == 74) || (y == 55 && x == 74) || (y == 56 && x == 74) || (y == 57 && x == 74) || (y == 58 && x == 74) || (y == 59 && x == 74) || (y == 60 && x == 74) || (y == 61 && x == 74) || (y == 62 && x == 74) || (y == 63 && x == 74) || (y == 0 && x == 75) || (y == 1 && x == 75) || (y == 2 && x == 75) || (y == 3 && x == 75) || (y == 4 && x == 75) || (y == 5 && x == 75) || (y == 6 && x == 75) || (y == 7 && x == 75) || (y == 8 && x == 75) || (y == 9 && x == 75) || (y == 10 && x == 75) || (y == 11 && x == 75) || (y == 12 && x == 75) || (y == 13 && x == 75) || (y == 14 && x == 75) || (y == 15 && x == 75) || (y == 16 && x == 75) || (y == 17 && x == 75) || (y == 18 && x == 75) || (y == 19 && x == 75) || (y == 20 && x == 75) || (y == 21 && x == 75) || (y == 22 && x == 75) || (y == 23 && x == 75) || (y == 24 && x == 75) || (y == 25 && x == 75) || (y == 26 && x == 75) || (y == 27 && x == 75) || (y == 28 && x == 75) || (y == 29 && x == 75) || (y == 30 && x == 75) || (y == 31 && x == 75) || (y == 32 && x == 75) || (y == 33 && x == 75) || (y == 34 && x == 75) || (y == 35 && x == 75) || (y == 36 && x == 75) || (y == 37 && x == 75) || (y == 38 && x == 75) || (y == 39 && x == 75) || (y == 40 && x == 75) || (y == 41 && x == 75) || (y == 42 && x == 75) || (y == 43 && x == 75) || (y == 44 && x == 75) || (y == 45 && x == 75) || (y == 46 && x == 75) || (y == 47 && x == 75) || (y == 48 && x == 75) || (y == 49 && x == 75) || (y == 50 && x == 75) || (y == 51 && x == 75) || (y == 52 && x == 75) || (y == 53 && x == 75) || (y == 54 && x == 75) || (y == 55 && x == 75) || (y == 56 && x == 75) || (y == 57 && x == 75) || (y == 58 && x == 75) || (y == 59 && x == 75) || (y == 60 && x == 75) || (y == 61 && x == 75) || (y == 62 && x == 75) || (y == 63 && x == 75) || (y == 0 && x == 76) || (y == 1 && x == 76) || (y == 2 && x == 76) || (y == 3 && x == 76) || (y == 4 && x == 76) || (y == 5 && x == 76) || (y == 6 && x == 76) || (y == 7 && x == 76) || (y == 8 && x == 76) || (y == 9 && x == 76) || (y == 10 && x == 76) || (y == 11 && x == 76) || (y == 12 && x == 76) || (y == 13 && x == 76) || (y == 14 && x == 76) || (y == 15 && x == 76) || (y == 16 && x == 76) || (y == 17 && x == 76) || (y == 18 && x == 76) || (y == 19 && x == 76) || (y == 20 && x == 76) || (y == 21 && x == 76) || (y == 22 && x == 76) || (y == 23 && x == 76) || (y == 24 && x == 76) || (y == 25 && x == 76) || (y == 26 && x == 76) || (y == 27 && x == 76) || (y == 28 && x == 76) || (y == 29 && x == 76) || (y == 30 && x == 76) || (y == 31 && x == 76) || (y == 32 && x == 76) || (y == 33 && x == 76) || (y == 34 && x == 76) || (y == 35 && x == 76) || (y == 36 && x == 76) || (y == 37 && x == 76) || (y == 38 && x == 76) || (y == 39 && x == 76) || (y == 40 && x == 76) || (y == 41 && x == 76) || (y == 42 && x == 76) || (y == 43 && x == 76) || (y == 44 && x == 76) || (y == 45 && x == 76) || (y == 46 && x == 76) || (y == 47 && x == 76) || (y == 48 && x == 76) || (y == 49 && x == 76) || (y == 50 && x == 76) || (y == 51 && x == 76) || (y == 52 && x == 76) || (y == 53 && x == 76) || (y == 54 && x == 76) || (y == 55 && x == 76) || (y == 56 && x == 76) || (y == 57 && x == 76) || (y == 58 && x == 76) || (y == 59 && x == 76) || (y == 60 && x == 76) || (y == 61 && x == 76) || (y == 62 && x == 76) || (y == 63 && x == 76) || (y == 0 && x == 77) || (y == 1 && x == 77) || (y == 2 && x == 77) || (y == 3 && x == 77) || (y == 4 && x == 77) || (y == 5 && x == 77) || (y == 6 && x == 77) || (y == 7 && x == 77) || (y == 8 && x == 77) || (y == 9 && x == 77) || (y == 10 && x == 77) || (y == 11 && x == 77) || (y == 12 && x == 77) || (y == 13 && x == 77) || (y == 14 && x == 77) || (y == 15 && x == 77) || (y == 16 && x == 77) || (y == 17 && x == 77) || (y == 18 && x == 77) || (y == 19 && x == 77) || (y == 20 && x == 77) || (y == 21 && x == 77) || (y == 22 && x == 77) || (y == 23 && x == 77) || (y == 24 && x == 77) || (y == 25 && x == 77) || (y == 26 && x == 77) || (y == 27 && x == 77) || (y == 28 && x == 77) || (y == 29 && x == 77) || (y == 30 && x == 77) || (y == 31 && x == 77) || (y == 32 && x == 77) || (y == 33 && x == 77) || (y == 34 && x == 77) || (y == 35 && x == 77) || (y == 36 && x == 77) || (y == 37 && x == 77) || (y == 38 && x == 77) || (y == 39 && x == 77) || (y == 40 && x == 77) || (y == 41 && x == 77) || (y == 42 && x == 77) || (y == 43 && x == 77) || (y == 44 && x == 77) || (y == 45 && x == 77) || (y == 46 && x == 77) || (y == 47 && x == 77) || (y == 48 && x == 77) || (y == 49 && x == 77) || (y == 50 && x == 77) || (y == 51 && x == 77) || (y == 52 && x == 77) || (y == 53 && x == 77) || (y == 54 && x == 77) || (y == 55 && x == 77) || (y == 56 && x == 77) || (y == 57 && x == 77) || (y == 58 && x == 77) || (y == 59 && x == 77) || (y == 60 && x == 77) || (y == 61 && x == 77) || (y == 62 && x == 77) || (y == 63 && x == 77) || (y == 0 && x == 78) || (y == 1 && x == 78) || (y == 2 && x == 78) || (y == 3 && x == 78) || (y == 4 && x == 78) || (y == 5 && x == 78) || (y == 6 && x == 78) || (y == 7 && x == 78) || (y == 8 && x == 78) || (y == 9 && x == 78) || (y == 10 && x == 78) || (y == 11 && x == 78) || (y == 12 && x == 78) || (y == 13 && x == 78) || (y == 14 && x == 78) || (y == 15 && x == 78) || (y == 16 && x == 78) || (y == 17 && x == 78) || (y == 18 && x == 78) || (y == 19 && x == 78) || (y == 20 && x == 78) || (y == 21 && x == 78) || (y == 22 && x == 78) || (y == 23 && x == 78) || (y == 24 && x == 78) || (y == 25 && x == 78) || (y == 26 && x == 78) || (y == 27 && x == 78) || (y == 28 && x == 78) || (y == 29 && x == 78) || (y == 30 && x == 78) || (y == 31 && x == 78) || (y == 32 && x == 78) || (y == 33 && x == 78) || (y == 34 && x == 78) || (y == 35 && x == 78) || (y == 36 && x == 78) || (y == 37 && x == 78) || (y == 38 && x == 78) || (y == 39 && x == 78) || (y == 40 && x == 78) || (y == 41 && x == 78) || (y == 42 && x == 78) || (y == 43 && x == 78) || (y == 44 && x == 78) || (y == 45 && x == 78) || (y == 46 && x == 78) || (y == 47 && x == 78) || (y == 48 && x == 78) || (y == 49 && x == 78) || (y == 50 && x == 78) || (y == 51 && x == 78) || (y == 52 && x == 78) || (y == 53 && x == 78) || (y == 54 && x == 78) || (y == 55 && x == 78) || (y == 56 && x == 78) || (y == 57 && x == 78) || (y == 58 && x == 78) || (y == 59 && x == 78) || (y == 60 && x == 78) || (y == 61 && x == 78) || (y == 62 && x == 78) || (y == 63 && x == 78) || (y == 0 && x == 79) || (y == 1 && x == 79) || (y == 2 && x == 79) || (y == 3 && x == 79) || (y == 4 && x == 79) || (y == 5 && x == 79) || (y == 6 && x == 79) || (y == 7 && x == 79) || (y == 8 && x == 79) || (y == 9 && x == 79) || (y == 10 && x == 79) || (y == 11 && x == 79) || (y == 12 && x == 79) || (y == 13 && x == 79) || (y == 14 && x == 79) || (y == 15 && x == 79) || (y == 16 && x == 79) || (y == 17 && x == 79) || (y == 18 && x == 79) || (y == 19 && x == 79) || (y == 20 && x == 79) || (y == 21 && x == 79) || (y == 22 && x == 79) || (y == 23 && x == 79) || (y == 24 && x == 79) || (y == 25 && x == 79) || (y == 26 && x == 79) || (y == 27 && x == 79) || (y == 28 && x == 79) || (y == 29 && x == 79) || (y == 30 && x == 79) || (y == 31 && x == 79) || (y == 32 && x == 79) || (y == 33 && x == 79) || (y == 34 && x == 79) || (y == 35 && x == 79) || (y == 36 && x == 79) || (y == 37 && x == 79) || (y == 38 && x == 79) || (y == 39 && x == 79) || (y == 40 && x == 79) || (y == 41 && x == 79) || (y == 42 && x == 79) || (y == 43 && x == 79) || (y == 44 && x == 79) || (y == 45 && x == 79) || (y == 46 && x == 79) || (y == 47 && x == 79) || (y == 48 && x == 79) || (y == 49 && x == 79) || (y == 50 && x == 79) || (y == 51 && x == 79) || (y == 52 && x == 79) || (y == 53 && x == 79) || (y == 54 && x == 79) || (y == 55 && x == 79) || (y == 56 && x == 79) || (y == 57 && x == 79) || (y == 58 && x == 79) || (y == 59 && x == 79) || (y == 60 && x == 79) || (y == 61 && x == 79) || (y == 62 && x == 79) || (y == 63 && x == 79) || (y == 0 && x == 80) || (y == 1 && x == 80) || (y == 2 && x == 80) || (y == 3 && x == 80) || (y == 4 && x == 80) || (y == 5 && x == 80) || (y == 6 && x == 80) || (y == 7 && x == 80) || (y == 8 && x == 80) || (y == 9 && x == 80) || (y == 10 && x == 80) || (y == 11 && x == 80) || (y == 12 && x == 80) || (y == 13 && x == 80) || (y == 14 && x == 80) || (y == 15 && x == 80) || (y == 16 && x == 80) || (y == 17 && x == 80) || (y == 18 && x == 80) || (y == 19 && x == 80) || (y == 20 && x == 80) || (y == 21 && x == 80) || (y == 22 && x == 80) || (y == 23 && x == 80) || (y == 24 && x == 80) || (y == 25 && x == 80) || (y == 26 && x == 80) || (y == 27 && x == 80) || (y == 28 && x == 80) || (y == 29 && x == 80) || (y == 30 && x == 80) || (y == 31 && x == 80) || (y == 32 && x == 80) || (y == 33 && x == 80) || (y == 34 && x == 80) || (y == 35 && x == 80) || (y == 36 && x == 80) || (y == 37 && x == 80) || (y == 38 && x == 80) || (y == 39 && x == 80) || (y == 40 && x == 80) || (y == 41 && x == 80) || (y == 42 && x == 80) || (y == 43 && x == 80) || (y == 44 && x == 80) || (y == 45 && x == 80) || (y == 46 && x == 80) || (y == 47 && x == 80) || (y == 48 && x == 80) || (y == 49 && x == 80) || (y == 50 && x == 80) || (y == 51 && x == 80) || (y == 52 && x == 80) || (y == 53 && x == 80) || (y == 54 && x == 80) || (y == 55 && x == 80) || (y == 56 && x == 80) || (y == 57 && x == 80) || (y == 58 && x == 80) || (y == 59 && x == 80) || (y == 60 && x == 80) || (y == 61 && x == 80) || (y == 62 && x == 80) || (y == 63 && x == 80) || (y == 0 && x == 81) || (y == 1 && x == 81) || (y == 2 && x == 81) || (y == 3 && x == 81) || (y == 4 && x == 81) || (y == 5 && x == 81) || (y == 6 && x == 81) || (y == 7 && x == 81) || (y == 8 && x == 81) || (y == 9 && x == 81) || (y == 10 && x == 81) || (y == 11 && x == 81) || (y == 12 && x == 81) || (y == 13 && x == 81) || (y == 14 && x == 81) || (y == 15 && x == 81) || (y == 16 && x == 81) || (y == 17 && x == 81) || (y == 18 && x == 81) || (y == 19 && x == 81) || (y == 20 && x == 81) || (y == 21 && x == 81) || (y == 22 && x == 81) || (y == 23 && x == 81) || (y == 24 && x == 81) || (y == 25 && x == 81) || (y == 26 && x == 81) || (y == 27 && x == 81) || (y == 28 && x == 81) || (y == 29 && x == 81) || (y == 30 && x == 81) || (y == 31 && x == 81) || (y == 32 && x == 81) || (y == 33 && x == 81) || (y == 34 && x == 81) || (y == 35 && x == 81) || (y == 36 && x == 81) || (y == 37 && x == 81) || (y == 38 && x == 81) || (y == 39 && x == 81) || (y == 40 && x == 81) || (y == 41 && x == 81) || (y == 42 && x == 81) || (y == 43 && x == 81) || (y == 44 && x == 81) || (y == 45 && x == 81) || (y == 46 && x == 81) || (y == 47 && x == 81) || (y == 48 && x == 81) || (y == 49 && x == 81) || (y == 50 && x == 81) || (y == 51 && x == 81) || (y == 52 && x == 81) || (y == 53 && x == 81) || (y == 54 && x == 81) || (y == 55 && x == 81) || (y == 56 && x == 81) || (y == 57 && x == 81) || (y == 58 && x == 81) || (y == 59 && x == 81) || (y == 60 && x == 81) || (y == 61 && x == 81) || (y == 62 && x == 81) || (y == 63 && x == 81) || (y == 0 && x == 82) || (y == 1 && x == 82) || (y == 2 && x == 82) || (y == 3 && x == 82) || (y == 4 && x == 82) || (y == 5 && x == 82) || (y == 6 && x == 82) || (y == 7 && x == 82) || (y == 8 && x == 82) || (y == 9 && x == 82) || (y == 10 && x == 82) || (y == 11 && x == 82) || (y == 12 && x == 82) || (y == 13 && x == 82) || (y == 14 && x == 82) || (y == 15 && x == 82) || (y == 16 && x == 82) || (y == 17 && x == 82) || (y == 18 && x == 82) || (y == 19 && x == 82) || (y == 20 && x == 82) || (y == 21 && x == 82) || (y == 22 && x == 82) || (y == 23 && x == 82) || (y == 24 && x == 82) || (y == 25 && x == 82) || (y == 26 && x == 82) || (y == 27 && x == 82) || (y == 28 && x == 82) || (y == 29 && x == 82) || (y == 30 && x == 82) || (y == 31 && x == 82) || (y == 32 && x == 82) || (y == 33 && x == 82) || (y == 34 && x == 82) || (y == 35 && x == 82) || (y == 36 && x == 82) || (y == 37 && x == 82) || (y == 38 && x == 82) || (y == 39 && x == 82) || (y == 40 && x == 82) || (y == 41 && x == 82) || (y == 42 && x == 82) || (y == 43 && x == 82) || (y == 44 && x == 82) || (y == 45 && x == 82) || (y == 46 && x == 82) || (y == 47 && x == 82) || (y == 48 && x == 82) || (y == 49 && x == 82) || (y == 50 && x == 82) || (y == 51 && x == 82) || (y == 52 && x == 82) || (y == 53 && x == 82) || (y == 54 && x == 82) || (y == 55 && x == 82) || (y == 56 && x == 82) || (y == 57 && x == 82) || (y == 58 && x == 82) || (y == 59 && x == 82) || (y == 60 && x == 82) || (y == 61 && x == 82) || (y == 62 && x == 82) || (y == 63 && x == 82) || (y == 0 && x == 83) || (y == 1 && x == 83) || (y == 2 && x == 83) || (y == 3 && x == 83) || (y == 4 && x == 83) || (y == 5 && x == 83) || (y == 6 && x == 83) || (y == 7 && x == 83) || (y == 8 && x == 83) || (y == 9 && x == 83) || (y == 10 && x == 83) || (y == 11 && x == 83) || (y == 12 && x == 83) || (y == 13 && x == 83) || (y == 14 && x == 83) || (y == 15 && x == 83) || (y == 16 && x == 83) || (y == 17 && x == 83) || (y == 18 && x == 83) || (y == 19 && x == 83) || (y == 20 && x == 83) || (y == 21 && x == 83) || (y == 22 && x == 83) || (y == 23 && x == 83) || (y == 24 && x == 83) || (y == 25 && x == 83) || (y == 26 && x == 83) || (y == 27 && x == 83) || (y == 28 && x == 83) || (y == 29 && x == 83) || (y == 30 && x == 83) || (y == 31 && x == 83) || (y == 32 && x == 83) || (y == 33 && x == 83) || (y == 34 && x == 83) || (y == 35 && x == 83) || (y == 36 && x == 83) || (y == 37 && x == 83) || (y == 38 && x == 83) || (y == 39 && x == 83) || (y == 40 && x == 83) || (y == 41 && x == 83) || (y == 42 && x == 83) || (y == 43 && x == 83) || (y == 44 && x == 83) || (y == 45 && x == 83) || (y == 46 && x == 83) || (y == 47 && x == 83) || (y == 48 && x == 83) || (y == 49 && x == 83) || (y == 50 && x == 83) || (y == 51 && x == 83) || (y == 52 && x == 83) || (y == 53 && x == 83) || (y == 54 && x == 83) || (y == 55 && x == 83) || (y == 56 && x == 83) || (y == 57 && x == 83) || (y == 58 && x == 83) || (y == 59 && x == 83) || (y == 60 && x == 83) || (y == 61 && x == 83) || (y == 62 && x == 83) || (y == 63 && x == 83) || (y == 0 && x == 84) || (y == 1 && x == 84) || (y == 2 && x == 84) || (y == 3 && x == 84) || (y == 4 && x == 84) || (y == 5 && x == 84) || (y == 6 && x == 84) || (y == 7 && x == 84) || (y == 8 && x == 84) || (y == 9 && x == 84) || (y == 10 && x == 84) || (y == 11 && x == 84) || (y == 12 && x == 84) || (y == 13 && x == 84) || (y == 14 && x == 84) || (y == 15 && x == 84) || (y == 16 && x == 84) || (y == 17 && x == 84) || (y == 18 && x == 84) || (y == 19 && x == 84) || (y == 20 && x == 84) || (y == 21 && x == 84) || (y == 22 && x == 84) || (y == 23 && x == 84) || (y == 24 && x == 84) || (y == 25 && x == 84) || (y == 26 && x == 84) || (y == 27 && x == 84) || (y == 28 && x == 84) || (y == 29 && x == 84) || (y == 30 && x == 84) || (y == 31 && x == 84) || (y == 32 && x == 84) || (y == 33 && x == 84) || (y == 34 && x == 84) || (y == 35 && x == 84) || (y == 36 && x == 84) || (y == 37 && x == 84) || (y == 38 && x == 84) || (y == 39 && x == 84) || (y == 40 && x == 84) || (y == 41 && x == 84) || (y == 42 && x == 84) || (y == 43 && x == 84) || (y == 44 && x == 84) || (y == 45 && x == 84) || (y == 46 && x == 84) || (y == 47 && x == 84) || (y == 48 && x == 84) || (y == 49 && x == 84) || (y == 50 && x == 84) || (y == 51 && x == 84) || (y == 52 && x == 84) || (y == 53 && x == 84) || (y == 54 && x == 84) || (y == 55 && x == 84) || (y == 56 && x == 84) || (y == 57 && x == 84) || (y == 58 && x == 84) || (y == 59 && x == 84) || (y == 60 && x == 84) || (y == 61 && x == 84) || (y == 62 && x == 84) || (y == 63 && x == 84) || (y == 0 && x == 85) || (y == 1 && x == 85) || (y == 2 && x == 85) || (y == 3 && x == 85) || (y == 4 && x == 85) || (y == 5 && x == 85) || (y == 6 && x == 85) || (y == 7 && x == 85) || (y == 8 && x == 85) || (y == 9 && x == 85) || (y == 10 && x == 85) || (y == 11 && x == 85) || (y == 12 && x == 85) || (y == 13 && x == 85) || (y == 14 && x == 85) || (y == 15 && x == 85) || (y == 16 && x == 85) || (y == 17 && x == 85) || (y == 18 && x == 85) || (y == 19 && x == 85) || (y == 20 && x == 85) || (y == 21 && x == 85) || (y == 22 && x == 85) || (y == 23 && x == 85) || (y == 24 && x == 85) || (y == 25 && x == 85) || (y == 26 && x == 85) || (y == 27 && x == 85) || (y == 28 && x == 85) || (y == 29 && x == 85) || (y == 30 && x == 85) || (y == 31 && x == 85) || (y == 32 && x == 85) || (y == 33 && x == 85) || (y == 34 && x == 85) || (y == 35 && x == 85) || (y == 36 && x == 85) || (y == 37 && x == 85) || (y == 38 && x == 85) || (y == 39 && x == 85) || (y == 40 && x == 85) || (y == 41 && x == 85) || (y == 42 && x == 85) || (y == 43 && x == 85) || (y == 44 && x == 85) || (y == 45 && x == 85) || (y == 46 && x == 85) || (y == 47 && x == 85) || (y == 48 && x == 85) || (y == 49 && x == 85) || (y == 50 && x == 85) || (y == 51 && x == 85) || (y == 52 && x == 85) || (y == 53 && x == 85) || (y == 54 && x == 85) || (y == 55 && x == 85) || (y == 56 && x == 85) || (y == 57 && x == 85) || (y == 58 && x == 85) || (y == 59 && x == 85) || (y == 60 && x == 85) || (y == 61 && x == 85) || (y == 62 && x == 85) || (y == 63 && x == 85) || (y == 0 && x == 86) || (y == 1 && x == 86) || (y == 2 && x == 86) || (y == 3 && x == 86) || (y == 4 && x == 86) || (y == 5 && x == 86) || (y == 6 && x == 86) || (y == 7 && x == 86) || (y == 8 && x == 86) || (y == 9 && x == 86) || (y == 10 && x == 86) || (y == 11 && x == 86) || (y == 12 && x == 86) || (y == 13 && x == 86) || (y == 14 && x == 86) || (y == 15 && x == 86) || (y == 16 && x == 86) || (y == 17 && x == 86) || (y == 18 && x == 86) || (y == 19 && x == 86) || (y == 20 && x == 86) || (y == 21 && x == 86) || (y == 22 && x == 86) || (y == 23 && x == 86) || (y == 24 && x == 86) || (y == 25 && x == 86) || (y == 26 && x == 86) || (y == 27 && x == 86) || (y == 28 && x == 86) || (y == 29 && x == 86) || (y == 30 && x == 86) || (y == 31 && x == 86) || (y == 32 && x == 86) || (y == 33 && x == 86) || (y == 34 && x == 86) || (y == 35 && x == 86) || (y == 36 && x == 86) || (y == 37 && x == 86) || (y == 38 && x == 86) || (y == 39 && x == 86) || (y == 40 && x == 86) || (y == 41 && x == 86) || (y == 42 && x == 86) || (y == 43 && x == 86) || (y == 44 && x == 86) || (y == 45 && x == 86) || (y == 46 && x == 86) || (y == 47 && x == 86) || (y == 48 && x == 86) || (y == 49 && x == 86) || (y == 50 && x == 86) || (y == 51 && x == 86) || (y == 52 && x == 86) || (y == 53 && x == 86) || (y == 54 && x == 86) || (y == 55 && x == 86) || (y == 56 && x == 86) || (y == 57 && x == 86) || (y == 58 && x == 86) || (y == 59 && x == 86) || (y == 60 && x == 86) || (y == 61 && x == 86) || (y == 62 && x == 86) || (y == 63 && x == 86) || (y == 0 && x == 87) || (y == 1 && x == 87) || (y == 2 && x == 87) || (y == 3 && x == 87) || (y == 4 && x == 87) || (y == 5 && x == 87) || (y == 6 && x == 87) || (y == 7 && x == 87) || (y == 8 && x == 87) || (y == 9 && x == 87) || (y == 10 && x == 87) || (y == 11 && x == 87) || (y == 12 && x == 87) || (y == 13 && x == 87) || (y == 14 && x == 87) || (y == 15 && x == 87) || (y == 16 && x == 87) || (y == 17 && x == 87) || (y == 18 && x == 87) || (y == 19 && x == 87) || (y == 20 && x == 87) || (y == 21 && x == 87) || (y == 22 && x == 87) || (y == 23 && x == 87) || (y == 24 && x == 87) || (y == 25 && x == 87) || (y == 26 && x == 87) || (y == 27 && x == 87) || (y == 28 && x == 87) || (y == 29 && x == 87) || (y == 30 && x == 87) || (y == 31 && x == 87) || (y == 32 && x == 87) || (y == 33 && x == 87) || (y == 34 && x == 87) || (y == 35 && x == 87) || (y == 36 && x == 87) || (y == 37 && x == 87) || (y == 38 && x == 87) || (y == 39 && x == 87) || (y == 40 && x == 87) || (y == 41 && x == 87) || (y == 42 && x == 87) || (y == 43 && x == 87) || (y == 44 && x == 87) || (y == 45 && x == 87) || (y == 46 && x == 87) || (y == 47 && x == 87) || (y == 48 && x == 87) || (y == 49 && x == 87) || (y == 50 && x == 87) || (y == 51 && x == 87) || (y == 52 && x == 87) || (y == 53 && x == 87) || (y == 54 && x == 87) || (y == 55 && x == 87) || (y == 56 && x == 87) || (y == 57 && x == 87) || (y == 58 && x == 87) || (y == 59 && x == 87) || (y == 60 && x == 87) || (y == 61 && x == 87) || (y == 62 && x == 87) || (y == 63 && x == 87) || (y == 0 && x == 88) || (y == 1 && x == 88) || (y == 2 && x == 88) || (y == 3 && x == 88) || (y == 4 && x == 88) || (y == 5 && x == 88) || (y == 6 && x == 88) || (y == 7 && x == 88) || (y == 8 && x == 88) || (y == 9 && x == 88) || (y == 10 && x == 88) || (y == 11 && x == 88) || (y == 12 && x == 88) || (y == 13 && x == 88) || (y == 14 && x == 88) || (y == 15 && x == 88) || (y == 16 && x == 88) || (y == 17 && x == 88) || (y == 18 && x == 88) || (y == 19 && x == 88) || (y == 20 && x == 88) || (y == 21 && x == 88) || (y == 22 && x == 88) || (y == 23 && x == 88) || (y == 24 && x == 88) || (y == 25 && x == 88) || (y == 26 && x == 88) || (y == 27 && x == 88) || (y == 28 && x == 88) || (y == 29 && x == 88) || (y == 30 && x == 88) || (y == 31 && x == 88) || (y == 32 && x == 88) || (y == 33 && x == 88) || (y == 34 && x == 88) || (y == 35 && x == 88) || (y == 36 && x == 88) || (y == 37 && x == 88) || (y == 38 && x == 88) || (y == 39 && x == 88) || (y == 40 && x == 88) || (y == 41 && x == 88) || (y == 42 && x == 88) || (y == 43 && x == 88) || (y == 44 && x == 88) || (y == 45 && x == 88) || (y == 46 && x == 88) || (y == 47 && x == 88) || (y == 48 && x == 88) || (y == 49 && x == 88) || (y == 50 && x == 88) || (y == 51 && x == 88) || (y == 52 && x == 88) || (y == 53 && x == 88) || (y == 54 && x == 88) || (y == 55 && x == 88) || (y == 56 && x == 88) || (y == 57 && x == 88) || (y == 58 && x == 88) || (y == 59 && x == 88) || (y == 60 && x == 88) || (y == 61 && x == 88) || (y == 62 && x == 88) || (y == 63 && x == 88) || (y == 0 && x == 89) || (y == 1 && x == 89) || (y == 2 && x == 89) || (y == 3 && x == 89) || (y == 4 && x == 89) || (y == 5 && x == 89) || (y == 6 && x == 89) || (y == 7 && x == 89) || (y == 8 && x == 89) || (y == 9 && x == 89) || (y == 10 && x == 89) || (y == 11 && x == 89) || (y == 12 && x == 89) || (y == 13 && x == 89) || (y == 14 && x == 89) || (y == 15 && x == 89) || (y == 16 && x == 89) || (y == 17 && x == 89) || (y == 18 && x == 89) || (y == 19 && x == 89) || (y == 20 && x == 89) || (y == 21 && x == 89) || (y == 22 && x == 89) || (y == 23 && x == 89) || (y == 24 && x == 89) || (y == 25 && x == 89) || (y == 26 && x == 89) || (y == 27 && x == 89) || (y == 28 && x == 89) || (y == 29 && x == 89) || (y == 30 && x == 89) || (y == 31 && x == 89) || (y == 32 && x == 89) || (y == 33 && x == 89) || (y == 34 && x == 89) || (y == 35 && x == 89) || (y == 36 && x == 89) || (y == 37 && x == 89) || (y == 38 && x == 89) || (y == 39 && x == 89) || (y == 40 && x == 89) || (y == 41 && x == 89) || (y == 42 && x == 89) || (y == 43 && x == 89) || (y == 44 && x == 89) || (y == 45 && x == 89) || (y == 46 && x == 89) || (y == 47 && x == 89) || (y == 48 && x == 89) || (y == 49 && x == 89) || (y == 50 && x == 89) || (y == 51 && x == 89) || (y == 52 && x == 89) || (y == 53 && x == 89) || (y == 54 && x == 89) || (y == 55 && x == 89) || (y == 56 && x == 89) || (y == 57 && x == 89) || (y == 58 && x == 89) || (y == 59 && x == 89) || (y == 60 && x == 89) || (y == 61 && x == 89) || (y == 62 && x == 89) || (y == 63 && x == 89) || (y == 0 && x == 90) || (y == 1 && x == 90) || (y == 2 && x == 90) || (y == 3 && x == 90) || (y == 4 && x == 90) || (y == 5 && x == 90) || (y == 6 && x == 90) || (y == 7 && x == 90) || (y == 8 && x == 90) || (y == 9 && x == 90) || (y == 10 && x == 90) || (y == 11 && x == 90) || (y == 12 && x == 90) || (y == 13 && x == 90) || (y == 14 && x == 90) || (y == 15 && x == 90) || (y == 16 && x == 90) || (y == 17 && x == 90) || (y == 18 && x == 90) || (y == 19 && x == 90) || (y == 20 && x == 90) || (y == 21 && x == 90) || (y == 22 && x == 90) || (y == 23 && x == 90) || (y == 24 && x == 90) || (y == 25 && x == 90) || (y == 26 && x == 90) || (y == 27 && x == 90) || (y == 28 && x == 90) || (y == 29 && x == 90) || (y == 30 && x == 90) || (y == 31 && x == 90) || (y == 32 && x == 90) || (y == 33 && x == 90) || (y == 34 && x == 90) || (y == 35 && x == 90) || (y == 36 && x == 90) || (y == 37 && x == 90) || (y == 38 && x == 90) || (y == 39 && x == 90) || (y == 40 && x == 90) || (y == 41 && x == 90) || (y == 42 && x == 90) || (y == 43 && x == 90) || (y == 44 && x == 90) || (y == 45 && x == 90) || (y == 46 && x == 90) || (y == 47 && x == 90) || (y == 48 && x == 90) || (y == 49 && x == 90) || (y == 50 && x == 90) || (y == 51 && x == 90) || (y == 52 && x == 90) || (y == 53 && x == 90) || (y == 54 && x == 90) || (y == 55 && x == 90) || (y == 56 && x == 90) || (y == 57 && x == 90) || (y == 58 && x == 90) || (y == 59 && x == 90) || (y == 60 && x == 90) || (y == 61 && x == 90) || (y == 62 && x == 90) || (y == 63 && x == 90) || (y == 0 && x == 91) || (y == 1 && x == 91) || (y == 2 && x == 91) || (y == 3 && x == 91) || (y == 4 && x == 91) || (y == 5 && x == 91) || (y == 6 && x == 91) || (y == 7 && x == 91) || (y == 8 && x == 91) || (y == 9 && x == 91) || (y == 10 && x == 91) || (y == 11 && x == 91) || (y == 12 && x == 91) || (y == 13 && x == 91) || (y == 14 && x == 91) || (y == 15 && x == 91) || (y == 16 && x == 91) || (y == 17 && x == 91) || (y == 18 && x == 91) || (y == 19 && x == 91) || (y == 20 && x == 91) || (y == 21 && x == 91) || (y == 22 && x == 91) || (y == 23 && x == 91) || (y == 24 && x == 91) || (y == 25 && x == 91) || (y == 26 && x == 91) || (y == 27 && x == 91) || (y == 28 && x == 91) || (y == 29 && x == 91) || (y == 30 && x == 91) || (y == 31 && x == 91) || (y == 32 && x == 91) || (y == 33 && x == 91) || (y == 34 && x == 91) || (y == 35 && x == 91) || (y == 36 && x == 91) || (y == 37 && x == 91) || (y == 38 && x == 91) || (y == 39 && x == 91) || (y == 40 && x == 91) || (y == 41 && x == 91) || (y == 42 && x == 91) || (y == 43 && x == 91) || (y == 44 && x == 91) || (y == 45 && x == 91) || (y == 46 && x == 91) || (y == 47 && x == 91) || (y == 48 && x == 91) || (y == 49 && x == 91) || (y == 50 && x == 91) || (y == 51 && x == 91) || (y == 52 && x == 91) || (y == 53 && x == 91) || (y == 54 && x == 91) || (y == 55 && x == 91) || (y == 56 && x == 91) || (y == 57 && x == 91) || (y == 58 && x == 91) || (y == 59 && x == 91) || (y == 60 && x == 91) || (y == 61 && x == 91) || (y == 62 && x == 91) || (y == 63 && x == 91) || (y == 0 && x == 92) || (y == 1 && x == 92) || (y == 2 && x == 92) || (y == 3 && x == 92) || (y == 4 && x == 92) || (y == 5 && x == 92) || (y == 6 && x == 92) || (y == 7 && x == 92) || (y == 8 && x == 92) || (y == 9 && x == 92) || (y == 10 && x == 92) || (y == 11 && x == 92) || (y == 12 && x == 92) || (y == 13 && x == 92) || (y == 14 && x == 92) || (y == 15 && x == 92) || (y == 16 && x == 92) || (y == 17 && x == 92) || (y == 18 && x == 92) || (y == 19 && x == 92) || (y == 20 && x == 92) || (y == 21 && x == 92) || (y == 22 && x == 92) || (y == 23 && x == 92) || (y == 24 && x == 92) || (y == 25 && x == 92) || (y == 26 && x == 92) || (y == 27 && x == 92) || (y == 28 && x == 92) || (y == 29 && x == 92) || (y == 30 && x == 92) || (y == 31 && x == 92) || (y == 32 && x == 92) || (y == 33 && x == 92) || (y == 34 && x == 92) || (y == 35 && x == 92) || (y == 36 && x == 92) || (y == 37 && x == 92) || (y == 38 && x == 92) || (y == 39 && x == 92) || (y == 40 && x == 92) || (y == 41 && x == 92) || (y == 42 && x == 92) || (y == 43 && x == 92) || (y == 44 && x == 92) || (y == 45 && x == 92) || (y == 46 && x == 92) || (y == 47 && x == 92) || (y == 48 && x == 92) || (y == 49 && x == 92) || (y == 50 && x == 92) || (y == 51 && x == 92) || (y == 52 && x == 92) || (y == 53 && x == 92) || (y == 54 && x == 92) || (y == 55 && x == 92) || (y == 56 && x == 92) || (y == 57 && x == 92) || (y == 58 && x == 92) || (y == 59 && x == 92) || (y == 60 && x == 92) || (y == 61 && x == 92) || (y == 62 && x == 92) || (y == 63 && x == 92) || (y == 0 && x == 93) || (y == 1 && x == 93) || (y == 2 && x == 93) || (y == 3 && x == 93) || (y == 4 && x == 93) || (y == 5 && x == 93) || (y == 6 && x == 93) || (y == 7 && x == 93) || (y == 8 && x == 93) || (y == 9 && x == 93) || (y == 10 && x == 93) || (y == 11 && x == 93) || (y == 12 && x == 93) || (y == 13 && x == 93) || (y == 14 && x == 93) || (y == 15 && x == 93) || (y == 16 && x == 93) || (y == 17 && x == 93) || (y == 18 && x == 93) || (y == 19 && x == 93) || (y == 20 && x == 93) || (y == 21 && x == 93) || (y == 22 && x == 93) || (y == 23 && x == 93) || (y == 24 && x == 93) || (y == 25 && x == 93) || (y == 26 && x == 93) || (y == 27 && x == 93) || (y == 28 && x == 93) || (y == 29 && x == 93) || (y == 30 && x == 93) || (y == 31 && x == 93) || (y == 32 && x == 93) || (y == 33 && x == 93) || (y == 34 && x == 93) || (y == 35 && x == 93) || (y == 36 && x == 93) || (y == 37 && x == 93) || (y == 38 && x == 93) || (y == 39 && x == 93) || (y == 40 && x == 93) || (y == 41 && x == 93) || (y == 42 && x == 93) || (y == 43 && x == 93) || (y == 44 && x == 93) || (y == 45 && x == 93) || (y == 46 && x == 93) || (y == 47 && x == 93) || (y == 48 && x == 93) || (y == 49 && x == 93) || (y == 50 && x == 93) || (y == 51 && x == 93) || (y == 52 && x == 93) || (y == 53 && x == 93) || (y == 54 && x == 93) || (y == 55 && x == 93) || (y == 56 && x == 93) || (y == 57 && x == 93) || (y == 58 && x == 93) || (y == 59 && x == 93) || (y == 60 && x == 93) || (y == 61 && x == 93) || (y == 62 && x == 93) || (y == 63 && x == 93) || (y == 0 && x == 94) || (y == 1 && x == 94) || (y == 2 && x == 94) || (y == 3 && x == 94) || (y == 4 && x == 94) || (y == 5 && x == 94) || (y == 6 && x == 94) || (y == 7 && x == 94) || (y == 8 && x == 94) || (y == 9 && x == 94) || (y == 10 && x == 94) || (y == 11 && x == 94) || (y == 12 && x == 94) || (y == 13 && x == 94) || (y == 14 && x == 94) || (y == 15 && x == 94) || (y == 16 && x == 94) || (y == 17 && x == 94) || (y == 18 && x == 94) || (y == 19 && x == 94) || (y == 20 && x == 94) || (y == 21 && x == 94) || (y == 22 && x == 94) || (y == 23 && x == 94) || (y == 24 && x == 94) || (y == 25 && x == 94) || (y == 26 && x == 94) || (y == 27 && x == 94) || (y == 28 && x == 94) || (y == 29 && x == 94) || (y == 30 && x == 94) || (y == 31 && x == 94) || (y == 32 && x == 94) || (y == 33 && x == 94) || (y == 34 && x == 94) || (y == 35 && x == 94) || (y == 36 && x == 94) || (y == 37 && x == 94) || (y == 38 && x == 94) || (y == 39 && x == 94) || (y == 40 && x == 94) || (y == 41 && x == 94) || (y == 42 && x == 94) || (y == 43 && x == 94) || (y == 44 && x == 94) || (y == 45 && x == 94) || (y == 46 && x == 94) || (y == 47 && x == 94) || (y == 48 && x == 94) || (y == 49 && x == 94) || (y == 50 && x == 94) || (y == 51 && x == 94) || (y == 52 && x == 94) || (y == 53 && x == 94) || (y == 54 && x == 94) || (y == 55 && x == 94) || (y == 56 && x == 94) || (y == 57 && x == 94) || (y == 58 && x == 94) || (y == 59 && x == 94) || (y == 60 && x == 94) || (y == 61 && x == 94) || (y == 62 && x == 94) || (y == 63 && x == 94) || (y == 0 && x == 95) || (y == 1 && x == 95) || (y == 2 && x == 95) || (y == 3 && x == 95) || (y == 4 && x == 95) || (y == 5 && x == 95) || (y == 6 && x == 95) || (y == 7 && x == 95) || (y == 8 && x == 95) || (y == 9 && x == 95) || (y == 10 && x == 95) || (y == 11 && x == 95) || (y == 12 && x == 95) || (y == 13 && x == 95) || (y == 14 && x == 95) || (y == 15 && x == 95) || (y == 16 && x == 95) || (y == 17 && x == 95) || (y == 18 && x == 95) || (y == 19 && x == 95) || (y == 20 && x == 95) || (y == 21 && x == 95) || (y == 22 && x == 95) || (y == 23 && x == 95) || (y == 24 && x == 95) || (y == 25 && x == 95) || (y == 26 && x == 95) || (y == 27 && x == 95) || (y == 28 && x == 95) || (y == 29 && x == 95) || (y == 30 && x == 95) || (y == 31 && x == 95) || (y == 32 && x == 95) || (y == 33 && x == 95) || (y == 34 && x == 95) || (y == 35 && x == 95) || (y == 36 && x == 95) || (y == 37 && x == 95) || (y == 38 && x == 95) || (y == 39 && x == 95) || (y == 40 && x == 95) || (y == 41 && x == 95) || (y == 42 && x == 95) || (y == 43 && x == 95) || (y == 44 && x == 95) || (y == 45 && x == 95) || (y == 46 && x == 95) || (y == 47 && x == 95) || (y == 48 && x == 95) || (y == 49 && x == 95) || (y == 50 && x == 95) || (y == 51 && x == 95) || (y == 52 && x == 95) || (y == 53 && x == 95) || (y == 54 && x == 95) || (y == 55 && x == 95) || (y == 56 && x == 95) || (y == 57 && x == 95) || (y == 58 && x == 95) || (y == 59 && x == 95) || (y == 60 && x == 95) || (y == 61 && x == 95) || (y == 62 && x == 95) || (y == 63 && x == 95)) oled_data <= 16'h29a6;
        else if ((y == 39 && x == 36)) oled_data <= 16'h265d;
        else if ((y == 23 && x == 35) || (y == 38 && x == 38) || (y == 36 && x == 41) || (y == 34 && x == 42) || (y == 36 && x == 42) || (y == 34 && x == 43) || (y == 36 && x == 43) || (y == 33 && x == 44) || (y == 34 && x == 44) || (y == 29 && x == 45) || (y == 32 && x == 45) || (y == 33 && x == 45) || (y == 29 && x == 46) || (y == 31 && x == 46) || (y == 32 && x == 46) || (y == 33 && x == 46) || (y == 30 && x == 47) || (y == 31 && x == 47) || (y == 30 && x == 48) || (y == 31 && x == 48) || (y == 30 && x == 49) || (y == 31 && x == 49) || (y == 30 && x == 50) || (y == 31 && x == 50) || (y == 34 && x == 50) || (y == 35 && x == 50) || (y == 30 && x == 51) || (y == 31 && x == 51) || (y == 32 && x == 51) || (y == 31 && x == 52) || (y == 32 && x == 52) || (y == 27 && x == 53) || (y == 32 && x == 53) || (y == 33 && x == 53) || (y == 34 && x == 53) || (y == 37 && x == 54) || (y == 40 && x == 57) || (y == 41 && x == 58) || (y == 43 && x == 59) || (y == 26 && x == 61) || (y == 39 && x == 61) || (y == 34 && x == 64)) oled_data <= 16'hf8a0;
        else if ((y == 34 && x == 63)) oled_data <= 16'h21cc;
        else if ((y == 45 && x == 30)) oled_data <= 16'h49eb;
        else if ((y == 45 && x == 39)) oled_data <= 16'hf300;
        else if ((y == 39 && x == 54) || (y == 38 && x == 55) || (y == 39 && x == 55) || (y == 34 && x == 57) || (y == 27 && x == 60)) oled_data <= 16'h980a;
        else if ((y == 46 && x == 60)) oled_data <= 16'h898e;
        else if ((y == 3 && x == 31) || (y == 4 && x == 31) || (y == 5 && x == 31) || (y == 6 && x == 31) || (y == 7 && x == 31) || (y == 8 && x == 31) || (y == 9 && x == 31) || (y == 10 && x == 31) || (y == 11 && x == 31) || (y == 12 && x == 31) || (y == 3 && x == 32) || (y == 4 && x == 32) || (y == 5 && x == 32) || (y == 6 && x == 32) || (y == 7 && x == 32) || (y == 8 && x == 32) || (y == 9 && x == 32) || (y == 10 && x == 32) || (y == 11 && x == 32) || (y == 12 && x == 32) || (y == 11 && x == 33) || (y == 12 && x == 33) || (y == 11 && x == 34) || (y == 12 && x == 34) || (y == 11 && x == 35) || (y == 12 && x == 35) || (y == 11 && x == 36) || (y == 12 && x == 36) || (y == 41 && x == 36) || (y == 11 && x == 37) || (y == 12 && x == 37) || (y == 11 && x == 38) || (y == 12 && x == 38) || (y == 59 && x == 40) || (y == 60 && x == 40) || (y == 61 && x == 40) || (y == 62 && x == 40) || (y == 63 && x == 40) || (y == 3 && x == 41) || (y == 4 && x == 41) || (y == 5 && x == 41) || (y == 6 && x == 41) || (y == 7 && x == 41) || (y == 8 && x == 41) || (y == 9 && x == 41) || (y == 10 && x == 41) || (y == 11 && x == 41) || (y == 12 && x == 41) || (y == 35 && x == 41) || (y == 59 && x == 41) || (y == 61 && x == 41) || (y == 62 && x == 41) || (y == 3 && x == 42) || (y == 4 && x == 42) || (y == 5 && x == 42) || (y == 6 && x == 42) || (y == 7 && x == 42) || (y == 8 && x == 42) || (y == 9 && x == 42) || (y == 10 && x == 42) || (y == 11 && x == 42) || (y == 12 && x == 42) || (y == 35 && x == 42) || (y == 46 && x == 42) || (y == 47 && x == 42) || (y == 59 && x == 42) || (y == 60 && x == 42) || (y == 61 && x == 42) || (y == 63 && x == 42) || (y == 3 && x == 43) || (y == 4 && x == 43) || (y == 11 && x == 43) || (y == 12 && x == 43) || (y == 25 && x == 43) || (y == 35 && x == 43) || (y == 46 && x == 43) || (y == 47 && x == 43) || (y == 48 && x == 43) || (y == 49 && x == 43) || (y == 50 && x == 43) || (y == 3 && x == 44) || (y == 4 && x == 44) || (y == 11 && x == 44) || (y == 12 && x == 44) || (y == 25 && x == 44) || (y == 47 && x == 44) || (y == 48 && x == 44) || (y == 49 && x == 44) || (y == 50 && x == 44) || (y == 59 && x == 44) || (y == 60 && x == 44) || (y == 61 && x == 44) || (y == 62 && x == 44) || (y == 63 && x == 44) || (y == 3 && x == 45) || (y == 4 && x == 45) || (y == 11 && x == 45) || (y == 12 && x == 45) || (y == 47 && x == 45) || (y == 48 && x == 45) || (y == 49 && x == 45) || (y == 50 && x == 45) || (y == 51 && x == 45) || (y == 59 && x == 45) || (y == 61 && x == 45) || (y == 63 && x == 45) || (y == 3 && x == 46) || (y == 4 && x == 46) || (y == 11 && x == 46) || (y == 12 && x == 46) || (y == 41 && x == 46) || (y == 46 && x == 46) || (y == 47 && x == 46) || (y == 48 && x == 46) || (y == 49 && x == 46) || (y == 50 && x == 46) || (y == 59 && x == 46) || (y == 61 && x == 46) || (y == 63 && x == 46) || (y == 3 && x == 47) || (y == 4 && x == 47) || (y == 5 && x == 47) || (y == 6 && x == 47) || (y == 7 && x == 47) || (y == 8 && x == 47) || (y == 9 && x == 47) || (y == 10 && x == 47) || (y == 11 && x == 47) || (y == 12 && x == 47) || (y == 41 && x == 47) || (y == 44 && x == 47) || (y == 46 && x == 47) || (y == 47 && x == 47) || (y == 48 && x == 47) || (y == 49 && x == 47) || (y == 50 && x == 47) || (y == 51 && x == 47) || (y == 3 && x == 48) || (y == 4 && x == 48) || (y == 5 && x == 48) || (y == 6 && x == 48) || (y == 7 && x == 48) || (y == 8 && x == 48) || (y == 9 && x == 48) || (y == 10 && x == 48) || (y == 11 && x == 48) || (y == 12 && x == 48) || (y == 41 && x == 48) || (y == 43 && x == 48) || (y == 44 && x == 48) || (y == 45 && x == 48) || (y == 46 && x == 48) || (y == 47 && x == 48) || (y == 48 && x == 48) || (y == 49 && x == 48) || (y == 50 && x == 48) || (y == 51 && x == 48) || (y == 59 && x == 48) || (y == 60 && x == 48) || (y == 61 && x == 48) || (y == 63 && x == 48) || (y == 41 && x == 49) || (y == 42 && x == 49) || (y == 43 && x == 49) || (y == 44 && x == 49) || (y == 45 && x == 49) || (y == 46 && x == 49) || (y == 47 && x == 49) || (y == 48 && x == 49) || (y == 49 && x == 49) || (y == 50 && x == 49) || (y == 51 && x == 49) || (y == 59 && x == 49) || (y == 61 && x == 49) || (y == 63 && x == 49) || (y == 41 && x == 50) || (y == 42 && x == 50) || (y == 44 && x == 50) || (y == 45 && x == 50) || (y == 46 && x == 50) || (y == 47 && x == 50) || (y == 48 && x == 50) || (y == 59 && x == 50) || (y == 61 && x == 50) || (y == 62 && x == 50) || (y == 63 && x == 50) || (y == 3 && x == 51) || (y == 4 && x == 51) || (y == 5 && x == 51) || (y == 6 && x == 51) || (y == 7 && x == 51) || (y == 8 && x == 51) || (y == 11 && x == 51) || (y == 12 && x == 51) || (y == 42 && x == 51) || (y == 44 && x == 51) || (y == 45 && x == 51) || (y == 46 && x == 51) || (y == 47 && x == 51) || (y == 48 && x == 51) || (y == 49 && x == 51) || (y == 3 && x == 52) || (y == 4 && x == 52) || (y == 5 && x == 52) || (y == 6 && x == 52) || (y == 7 && x == 52) || (y == 8 && x == 52) || (y == 11 && x == 52) || (y == 12 && x == 52) || (y == 46 && x == 52) || (y == 47 && x == 52) || (y == 49 && x == 52) || (y == 59 && x == 52) || (y == 60 && x == 52) || (y == 61 && x == 52) || (y == 62 && x == 52) || (y == 63 && x == 52) || (y == 3 && x == 53) || (y == 4 && x == 53) || (y == 7 && x == 53) || (y == 8 && x == 53) || (y == 11 && x == 53) || (y == 12 && x == 53) || (y == 35 && x == 53) || (y == 59 && x == 53) || (y == 61 && x == 53) || (y == 63 && x == 53) || (y == 3 && x == 54) || (y == 4 && x == 54) || (y == 7 && x == 54) || (y == 8 && x == 54) || (y == 11 && x == 54) || (y == 12 && x == 54) || (y == 59 && x == 54) || (y == 61 && x == 54) || (y == 63 && x == 54) || (y == 3 && x == 55) || (y == 4 && x == 55) || (y == 7 && x == 55) || (y == 8 && x == 55) || (y == 11 && x == 55) || (y == 12 && x == 55) || (y == 3 && x == 56) || (y == 4 && x == 56) || (y == 7 && x == 56) || (y == 8 && x == 56) || (y == 11 && x == 56) || (y == 12 && x == 56) || (y == 59 && x == 56) || (y == 3 && x == 57) || (y == 4 && x == 57) || (y == 7 && x == 57) || (y == 8 && x == 57) || (y == 9 && x == 57) || (y == 10 && x == 57) || (y == 11 && x == 57) || (y == 12 && x == 57) || (y == 59 && x == 57) || (y == 60 && x == 57) || (y == 61 && x == 57) || (y == 62 && x == 57) || (y == 63 && x == 57) || (y == 3 && x == 58) || (y == 4 && x == 58) || (y == 7 && x == 58) || (y == 8 && x == 58) || (y == 9 && x == 58) || (y == 10 && x == 58) || (y == 11 && x == 58) || (y == 12 && x == 58) || (y == 59 && x == 58) || (y == 47 && x == 60) || (y == 3 && x == 61) || (y == 4 && x == 61) || (y == 5 && x == 61) || (y == 6 && x == 61) || (y == 7 && x == 61) || (y == 8 && x == 61) || (y == 9 && x == 61) || (y == 10 && x == 61) || (y == 11 && x == 61) || (y == 12 && x == 61) || (y == 47 && x == 61) || (y == 3 && x == 62) || (y == 4 && x == 62) || (y == 5 && x == 62) || (y == 6 && x == 62) || (y == 7 && x == 62) || (y == 8 && x == 62) || (y == 9 && x == 62) || (y == 10 && x == 62) || (y == 11 && x == 62) || (y == 12 && x == 62) || (y == 47 && x == 62) || (y == 3 && x == 63) || (y == 4 && x == 63) || (y == 7 && x == 63) || (y == 8 && x == 63) || (y == 11 && x == 63) || (y == 12 && x == 63) || (y == 3 && x == 64) || (y == 4 && x == 64) || (y == 7 && x == 64) || (y == 8 && x == 64) || (y == 11 && x == 64) || (y == 12 && x == 64) || (y == 3 && x == 65) || (y == 4 && x == 65) || (y == 7 && x == 65) || (y == 8 && x == 65) || (y == 11 && x == 65) || (y == 12 && x == 65) || (y == 3 && x == 66) || (y == 4 && x == 66) || (y == 7 && x == 66) || (y == 8 && x == 66) || (y == 11 && x == 66) || (y == 12 && x == 66) || (y == 3 && x == 67) || (y == 4 && x == 67) || (y == 7 && x == 67) || (y == 8 && x == 67) || (y == 11 && x == 67) || (y == 12 && x == 67) || (y == 3 && x == 68) || (y == 4 && x == 68) || (y == 7 && x == 68) || (y == 8 && x == 68) || (y == 11 && x == 68) || (y == 12 && x == 68)) oled_data <= 16'hffff;
        else if ((y == 28 && x == 38) || (y == 39 && x == 38) || (y == 29 && x == 48) || (y == 29 && x == 49) || (y == 29 && x == 50) || (y == 30 && x == 52)) oled_data <= 16'ha808;
        else if ((y == 37 && x == 45) || (y == 37 && x == 46) || (y == 37 && x == 47)) oled_data <= 16'hfc00;
        else if ((y == 33 && x == 52)) oled_data <= 16'he082;
        else if ((y == 34 && x == 38)) oled_data <= 16'h506c;
        else if ((y == 44 && x == 54)) oled_data <= 16'hda84;
        else if ((y == 36 && x == 51) || (y == 42 && x == 59) || (y == 33 && x == 64)) oled_data <= 16'hf8c0;
        else if ((y == 43 && x == 29) || (y == 25 && x == 31)) oled_data <= 16'h316b;
        else if ((y == 34 && x == 25)) oled_data <= 16'h31c6;
        else if ((y == 52 && x == 50) || (y == 49 && x == 58)) oled_data <= 16'hfa98;
        else if ((y == 42 && x == 27) || (y == 43 && x == 27) || (y == 44 && x == 27) || (y == 42 && x == 28) || (y == 43 && x == 28) || (y == 44 && x == 28) || (y == 32 && x == 29) || (y == 33 && x == 29) || (y == 34 && x == 29) || (y == 39 && x == 29) || (y == 29 && x == 30) || (y == 30 && x == 30) || (y == 31 && x == 30) || (y == 32 && x == 30) || (y == 33 && x == 30) || (y == 34 && x == 30) || (y == 38 && x == 30) || (y == 39 && x == 30) || (y == 40 && x == 30) || (y == 44 && x == 30) || (y == 28 && x == 31) || (y == 29 && x == 31) || (y == 30 && x == 31) || (y == 31 && x == 31) || (y == 32 && x == 31) || (y == 33 && x == 31) || (y == 34 && x == 31) || (y == 37 && x == 31) || (y == 38 && x == 31) || (y == 39 && x == 31) || (y == 40 && x == 31) || (y == 44 && x == 31) || (y == 45 && x == 31) || (y == 27 && x == 32) || (y == 28 && x == 32) || (y == 29 && x == 32) || (y == 30 && x == 32) || (y == 31 && x == 32) || (y == 32 && x == 32) || (y == 33 && x == 32) || (y == 34 && x == 32) || (y == 36 && x == 32) || (y == 37 && x == 32) || (y == 38 && x == 32) || (y == 39 && x == 32) || (y == 40 && x == 32) || (y == 41 && x == 32) || (y == 43 && x == 32) || (y == 26 && x == 33) || (y == 27 && x == 33) || (y == 28 && x == 33) || (y == 29 && x == 33) || (y == 30 && x == 33) || (y == 31 && x == 33) || (y == 32 && x == 33) || (y == 41 && x == 33) || (y == 25 && x == 34) || (y == 26 && x == 34) || (y == 27 && x == 34) || (y == 28 && x == 34) || (y == 29 && x == 34) || (y == 30 && x == 34) || (y == 31 && x == 34) || (y == 33 && x == 34) || (y == 34 && x == 34) || (y == 45 && x == 34) || (y == 25 && x == 35) || (y == 26 && x == 35) || (y == 27 && x == 35) || (y == 28 && x == 35) || (y == 29 && x == 35) || (y == 30 && x == 35) || (y == 31 && x == 35) || (y == 32 && x == 35) || (y == 33 && x == 35) || (y == 45 && x == 35) || (y == 46 && x == 35) || (y == 26 && x == 36) || (y == 27 && x == 36) || (y == 28 && x == 36) || (y == 29 && x == 36) || (y == 30 && x == 36) || (y == 31 && x == 36) || (y == 32 && x == 36) || (y == 34 && x == 36) || (y == 28 && x == 37) || (y == 30 && x == 37) || (y == 31 && x == 37) || (y == 24 && x == 38) || (y == 25 && x == 38) || (y == 26 && x == 38) || (y == 30 && x == 38) || (y == 31 && x == 38) || (y == 33 && x == 38) || (y == 24 && x == 39) || (y == 25 && x == 39) || (y == 26 && x == 39) || (y == 27 && x == 39) || (y == 28 && x == 39) || (y == 31 && x == 39) || (y == 24 && x == 40) || (y == 25 && x == 40) || (y == 26 && x == 40) || (y == 27 && x == 40) || (y == 28 && x == 40) || (y == 29 && x == 40) || (y == 23 && x == 41) || (y == 24 && x == 41) || (y == 25 && x == 41) || (y == 26 && x == 41) || (y == 27 && x == 41) || (y == 28 && x == 41) || (y == 29 && x == 41) || (y == 23 && x == 42) || (y == 24 && x == 42) || (y == 25 && x == 42) || (y == 22 && x == 43) || (y == 23 && x == 43) || (y == 24 && x == 43) || (y == 26 && x == 43) || (y == 22 && x == 44) || (y == 23 && x == 44) || (y == 24 && x == 44) || (y == 26 && x == 44) || (y == 22 && x == 45) || (y == 23 && x == 45) || (y == 24 && x == 45) || (y == 27 && x == 45) || (y == 21 && x == 46) || (y == 22 && x == 46) || (y == 23 && x == 46) || (y == 21 && x == 47) || (y == 22 && x == 47) || (y == 24 && x == 47) || (y == 21 && x == 48) || (y == 22 && x == 48) || (y == 22 && x == 49) || (y == 22 && x == 50) || (y == 22 && x == 51) || (y == 23 && x == 52) || (y == 24 && x == 52) || (y == 23 && x == 53) || (y == 24 && x == 53) || (y == 24 && x == 54) || (y == 25 && x == 54) || (y == 25 && x == 55) || (y == 28 && x == 55) || (y == 29 && x == 55) || (y == 30 && x == 55) || (y == 27 && x == 56) || (y == 29 && x == 56) || (y == 30 && x == 56) || (y == 31 && x == 56) || (y == 32 && x == 56) || (y == 31 && x == 57) || (y == 32 && x == 57) || (y == 33 && x == 57) || (y == 27 && x == 58) || (y == 28 && x == 58) || (y == 29 && x == 58) || (y == 30 && x == 58) || (y == 30 && x == 60) || (y == 32 && x == 60) || (y == 30 && x == 61) || (y == 31 && x == 62) || (y == 37 && x == 62) || (y == 38 && x == 62) || (y == 32 && x == 63) || (y == 33 && x == 63) || (y == 36 && x == 63) || (y == 37 && x == 63) || (y == 32 && x == 64) || (y == 36 && x == 64) || (y == 37 && x == 64) || (y == 38 && x == 64) || (y == 39 && x == 64) || (y == 40 && x == 64) || (y == 41 && x == 64) || (y == 36 && x == 65) || (y == 37 && x == 65) || (y == 38 && x == 65) || (y == 39 && x == 65) || (y == 40 && x == 65) || (y == 36 && x == 66) || (y == 37 && x == 66) || (y == 38 && x == 66) || (y == 39 && x == 66) || (y == 37 && x == 67) || (y == 38 && x == 67) || (y == 39 && x == 67) || (y == 38 && x == 68) || (y == 39 && x == 68)) oled_data <= 16'h29cb;
        else if ((y == 36 && x == 62)) oled_data <= 16'h8146;
        else if ((y == 38 && x == 35) || (y == 25 && x == 36) || (y == 36 && x == 36) || (y == 37 && x == 36) || (y == 38 && x == 36) || (y == 35 && x == 37) || (y == 36 && x == 37) || (y == 37 && x == 37) || (y == 38 && x == 37) || (y == 39 && x == 37) || (y == 40 && x == 37) || (y == 36 && x == 38) || (y == 37 && x == 38) || (y == 40 && x == 38) || (y == 35 && x == 39) || (y == 36 && x == 39) || (y == 39 && x == 39) || (y == 38 && x == 40) || (y == 37 && x == 41) || (y == 33 && x == 42) || (y == 29 && x == 43) || (y == 32 && x == 43) || (y == 33 && x == 43) || (y == 29 && x == 44) || (y == 31 && x == 44) || (y == 32 && x == 44) || (y == 28 && x == 45) || (y == 31 && x == 45) || (y == 28 && x == 47) || (y == 29 && x == 47) || (y == 25 && x == 48) || (y == 28 && x == 48) || (y == 25 && x == 49) || (y == 27 && x == 49) || (y == 28 && x == 49) || (y == 27 && x == 50) || (y == 28 && x == 50) || (y == 27 && x == 51) || (y == 28 && x == 51) || (y == 29 && x == 51) || (y == 28 && x == 52) || (y == 29 && x == 52) || (y == 34 && x == 52) || (y == 35 && x == 52) || (y == 30 && x == 53) || (y == 31 && x == 53) || (y == 28 && x == 54) || (y == 34 && x == 54) || (y == 36 && x == 54) || (y == 37 && x == 55) || (y == 40 && x == 55) || (y == 36 && x == 56) || (y == 37 && x == 56) || (y == 38 && x == 56) || (y == 39 && x == 56) || (y == 40 && x == 56) || (y == 41 && x == 56) || (y == 35 && x == 57) || (y == 39 && x == 57) || (y == 41 && x == 57) || (y == 42 && x == 57) || (y == 39 && x == 58) || (y == 40 && x == 58) || (y == 38 && x == 59) || (y == 39 && x == 59) || (y == 40 && x == 59) || (y == 41 && x == 59) || (y == 29 && x == 60) || (y == 39 && x == 60) || (y == 40 && x == 60) || (y == 41 && x == 60) || (y == 42 && x == 60) || (y == 25 && x == 61) || (y == 28 && x == 61) || (y == 41 && x == 61) || (y == 42 && x == 61) || (y == 34 && x == 65)) oled_data <= 16'ha009;
        else if ((y == 46 && x == 54)) oled_data <= 16'hfd80;
        else if ((y == 51 && x == 50)) oled_data <= 16'hff98;
        else if ((y == 46 && x == 63)) oled_data <= 16'ha9f0;
        else if ((y == 51 && x == 62)) oled_data <= 16'hc232;
        else if ((y == 25 && x == 45) || (y == 28 && x == 57)) oled_data <= 16'hf1f;
        else if ((y == 30 && x == 46)) oled_data <= 16'hc846;
        else if ((y == 47 && x == 59)) oled_data <= 16'h71f;
        else if ((y == 36 && x == 72) || (y == 38 && x == 73) || (y == 39 && x == 73) || (y == 40 && x == 73)) oled_data <= 16'h2910;
        else if ((y == 27 && x == 48)) oled_data <= 16'h48cd;
        else if ((y == 44 && x == 59)) oled_data <= 16'h7170;
        else if ((y == 26 && x == 56) || (y == 37 && x == 73)) oled_data <= 16'h296a;
        else if ((y == 26 && x == 60) || (y == 26 && x == 68)) oled_data <= 16'h3188;
        else if ((y == 45 && x == 62)) oled_data <= 16'h4477;
        else if ((y == 37 && x == 72)) oled_data <= 16'h28d1;
        else if ((y == 38 && x == 39) || (y == 32 && x == 41) || (y == 38 && x == 60)) oled_data <= 16'hc046;
        else if ((y == 45 && x == 25) || (y == 45 && x == 71)) oled_data <= 16'h28d4;
        else if ((y == 37 && x == 40)) oled_data <= 16'hf241;
        else if ((y == 40 && x == 42)) oled_data <= 16'hfe20;
        else if ((y == 46 && x == 30) || (y == 45 && x == 63)) oled_data <= 16'hf297;
        else if ((y == 45 && x == 53)) oled_data <= 16'ha3ea;
        else if ((y == 45 && x == 37) || (y == 46 && x == 37) || (y == 47 && x == 37) || (y == 45 && x == 38) || (y == 46 && x == 38) || (y == 47 && x == 38) || (y == 48 && x == 38) || (y == 41 && x == 39) || (y == 42 && x == 39) || (y == 43 && x == 39) || (y == 39 && x == 40) || (y == 40 && x == 40) || (y == 41 && x == 40) || (y == 42 && x == 40) || (y == 43 && x == 40) || (y == 38 && x == 41) || (y == 39 && x == 41) || (y == 40 && x == 41) || (y == 43 && x == 41) || (y == 38 && x == 42) || (y == 39 && x == 42) || (y == 42 && x == 42) || (y == 43 && x == 42) || (y == 37 && x == 43) || (y == 38 && x == 43) || (y == 39 && x == 43) || (y == 41 && x == 43) || (y == 42 && x == 43) || (y == 43 && x == 43) || (y == 37 && x == 44) || (y == 38 && x == 44) || (y == 41 && x == 44) || (y == 35 && x == 45) || (y == 36 && x == 45) || (y == 34 && x == 46) || (y == 35 && x == 46) || (y == 36 && x == 46) || (y == 32 && x == 47) || (y == 34 && x == 47) || (y == 35 && x == 47) || (y == 36 && x == 47) || (y == 32 && x == 48) || (y == 34 && x == 48) || (y == 35 && x == 48) || (y == 36 && x == 48) || (y == 37 && x == 48) || (y == 33 && x == 49) || (y == 34 && x == 49) || (y == 35 && x == 49) || (y == 36 && x == 49) || (y == 37 && x == 49) || (y == 39 && x == 49) || (y == 32 && x == 50) || (y == 36 && x == 50) || (y == 37 && x == 50) || (y == 39 && x == 50) || (y == 37 && x == 51) || (y == 40 && x == 51) || (y == 36 && x == 52) || (y == 37 && x == 52) || (y == 38 && x == 52) || (y == 39 && x == 52) || (y == 41 && x == 52) || (y == 37 && x == 53) || (y == 38 && x == 53) || (y == 39 && x == 53) || (y == 40 && x == 53) || (y == 41 && x == 53) || (y == 41 && x == 54) || (y == 42 && x == 54) || (y == 42 && x == 55) || (y == 43 && x == 55) || (y == 46 && x == 55) || (y == 42 && x == 56) || (y == 43 && x == 56) || (y == 46 && x == 56) || (y == 47 && x == 56) || (y == 48 && x == 56) || (y == 45 && x == 57) || (y == 46 && x == 57) || (y == 32 && x == 58) || (y == 42 && x == 58) || (y == 43 && x == 58) || (y == 28 && x == 60)) oled_data <= 16'hfb00;
        else if ((y == 19 && x == 39)) oled_data <= 16'h3169;
        else if ((y == 52 && x == 40) || (y == 52 && x == 41) || (y == 52 && x == 55) || (y == 52 && x == 60)) oled_data <= 16'h81ed;
        else if ((y == 49 && x == 34)) oled_data <= 16'h4a0b;
        else if ((y == 49 && x == 25) || (y == 46 && x == 26) || (y == 47 && x == 27) || (y == 57 && x == 40) || (y == 56 && x == 46) || (y == 15 && x == 50) || (y == 57 && x == 50) || (y == 57 && x == 51) || (y == 56 && x == 52) || (y == 54 && x == 61) || (y == 27 && x == 62) || (y == 24 && x == 67) || (y == 29 && x == 71) || (y == 30 && x == 72)) oled_data <= 16'h29a8;
        else if ((y == 46 && x == 27) || (y == 47 && x == 31) || (y == 46 && x == 67)) oled_data <= 16'h61ec;
        else if ((y == 32 && x == 39)) oled_data <= 16'h269e;
        else if ((y == 26 && x == 62)) oled_data <= 16'h58e8;
        else if ((y == 49 && x == 32) || (y == 46 && x == 33) || (y == 50 && x == 34) || (y == 48 && x == 59) || (y == 50 && x == 63)) oled_data <= 16'hfab9;
        else if ((y == 27 && x == 37) || (y == 28 && x == 59)) oled_data <= 16'h21eb;
        else if ((y == 48 && x == 33) || (y == 48 && x == 35) || (y == 48 && x == 36) || (y == 48 && x == 61)) oled_data <= 16'h91ad;
        else if ((y == 49 && x == 39) || (y == 49 && x == 62)) oled_data <= 16'h99cd;
        else if ((y == 30 && x == 41)) oled_data <= 16'hcdd;
        else if ((y == 38 && x == 51)) oled_data <= 16'hfc20;
        else if ((y == 40 && x == 39)) oled_data <= 16'hf8e0;
        else if ((y == 42 && x == 72)) oled_data <= 16'h4152;
        else if ((y == 46 && x == 23) || (y == 49 && x == 63) || (y == 52 && x == 65)) oled_data <= 16'h49ea;
        else if ((y == 24 && x == 36) || (y == 41 && x == 41) || (y == 44 && x == 41)) oled_data <= 16'hfd60;
        else if ((y == 44 && x == 56)) oled_data <= 16'h4994;
        else oled_data <= 16'hffff;
    end
endmodule
