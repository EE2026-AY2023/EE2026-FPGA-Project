`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 29.03.2023 23:07:20
// Design Name: 
// Module Name: ftb_start_screen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//bomb sprite credit: https://www.kindpng.com/imgv/iTJRhw_bomb-omb-pixel-art-hd-png-download/
//alphabets credits: https://www.alamy.com/stock-image-pixel-alphabet-isolated-digital-font-169448226.html?imageid=0C5C03FE-8B9C-4229-B30A-F896C25571CC&p=358500&pn=2&searchId=38fc8283011d9b09d3e1276b9e308ec5&searchtype=0

module ftb_start_screen(
    input clock,
    input [6:0] x, y,
    output reg [15:0] oled_data = 0
    );
    reg [31:0] count = 0;
    always @(posedge clock) begin
        if ((y == 55 && x == 43)) oled_data <= 16'h8c51;
        else if ((y == 43 && x == 13) || (y == 42 && x == 24)) oled_data <= 16'hde7a;
        else if ((y == 25 && x == 23)) oled_data <= 16'he6bb;
        else if ((y == 20 && x == 23) || (y == 21 && x == 23)) oled_data <= 16'hdeda;
        else if ((y == 11 && x == 18) || (y == 11 && x == 20)) oled_data <= 16'h9410;
        else if ((y == 37 && x == 5) || (y == 20 && x == 18) || (y == 21 && x == 18) || (y == 22 && x == 18) || (y == 29 && x == 18) || (y == 30 && x == 18) || (y == 37 && x == 35)) oled_data <= 16'h5249;
        else if ((y == 24 && x == 18) || (y == 28 && x == 18)) oled_data <= 16'h5229;
        else if ((y == 40 && x == 9) || (y == 43 && x == 9) || (y == 24 && x == 17) || (y == 38 && x == 26) || (y == 40 && x == 39) || (y == 43 && x == 39)) oled_data <= 16'h28e3;
        else if ((y == 39 && x == 26)) oled_data <= 16'h20c3;
        else if ((y == 15 && x == 33)) oled_data <= 16'hbdf7;
        else if ((y == 38 && x == 10) || (y == 38 && x == 40)) oled_data <= 16'h3144;
        else if ((y == 25 && x == 16)) oled_data <= 16'h1841;
        else if ((y == 20 && x == 7) || (y == 21 && x == 7) || (y == 22 && x == 7) || (y == 24 && x == 7) || (y == 29 && x == 7) || (y == 30 && x == 7) || (y == 30 && x == 24) || (y == 54 && x == 39) || (y == 55 && x == 39) || (y == 56 && x == 39) || (y == 59 && x == 39) || (y == 54 && x == 54) || (y == 55 && x == 54) || (y == 56 && x == 54) || (y == 59 && x == 54)) oled_data <= 16'h1041;
        else if ((y == 6 && x == 29)) oled_data <= 16'h39a5;
        else if ((y == 28 && x == 6)) oled_data <= 16'hce38;
        else if ((y == 24 && x == 23) || (y == 26 && x == 23) || (y == 27 && x == 23) || (y == 28 && x == 23)) oled_data <= 16'he6da;
        else if ((y == 26 && x == 14)) oled_data <= 16'hf79d;
        else if ((y == 8 && x == 5) || (y == 11 && x == 19) || (y == 27 && x == 19) || (y == 8 && x == 28) || (y == 9 && x == 28) || (y == 10 && x == 28) || (y == 11 && x == 28)) oled_data <= 16'h8c10;
        else if ((y == 6 && x == 28)) oled_data <= 16'h9492;
        else if ((y == 57 && x == 50)) oled_data <= 16'h9cb3;
        else if ((y == 21 && x == 6) || (y == 27 && x == 6)) oled_data <= 16'hce18;
        else if ((y == 14 && x == 4) || (y == 7 && x == 5) || (y == 11 && x == 13) || (y == 27 && x == 13) || (y == 11 && x == 14) || (y == 27 && x == 14) || (y == 43 && x == 14) || (y == 9 && x == 18) || (y == 9 && x == 19) || (y == 9 && x == 20) || (y == 9 && x == 22) || (y == 9 && x == 23) || (y == 21 && x == 24) || (y == 7 && x == 27) || (y == 41 && x == 30)) oled_data <= 16'h800;
        else if ((y == 22 && x == 5) || (y == 11 && x == 6) || (y == 43 && x == 6) || (y == 9 && x == 9) || (y == 22 && x == 9) || (y == 22 && x == 10) || (y == 31 && x == 13) || (y == 15 && x == 14) || (y == 31 && x == 14) || (y == 4 && x == 15) || (y == 12 && x == 15) || (y == 15 && x == 15) || (y == 21 && x == 15) || (y == 22 && x == 15) || (y == 23 && x == 15) || (y == 27 && x == 15) || (y == 28 && x == 15) || (y == 29 && x == 15) || (y == 30 && x == 15) || (y == 31 && x == 15) || (y == 31 && x == 18) || (y == 15 && x == 19) || (y == 31 && x == 19) || (y == 15 && x == 23) || (y == 9 && x == 24) || (y == 10 && x == 24) || (y == 15 && x == 24) || (y == 36 && x == 24) || (y == 47 && x == 24) || (y == 47 && x == 25) || (y == 40 && x == 26) || (y == 47 && x == 30) || (y == 55 && x == 34) || (y == 55 && x == 35) || (y == 43 && x == 36) || (y == 55 && x == 38) || (y == 55 && x == 40) || (y == 55 && x == 49) || (y == 55 && x == 53) || (y == 55 && x == 55)) oled_data <= 16'had75;
        else if ((y == 20 && x == 6)) oled_data <= 16'hd638;
        else if ((y == 45 && x == 9) || (y == 45 && x == 39)) oled_data <= 16'h2904;
        else if ((y == 39 && x == 24)) oled_data <= 16'h1840;
        else if ((y == 6 && x == 27)) oled_data <= 16'h41a7;
        else if ((y == 39 && x == 6) || (y == 40 && x == 6) || (y == 44 && x == 6) || (y == 11 && x == 7) || (y == 31 && x == 7) || (y == 43 && x == 7) || (y == 11 && x == 8) || (y == 31 && x == 8) || (y == 10 && x == 9) || (y == 11 && x == 9) || (y == 5 && x == 10) || (y == 6 && x == 10) || (y == 47 && x == 14) || (y == 20 && x == 15) || (y == 47 && x == 15) || (y == 38 && x == 16) || (y == 47 && x == 16) || (y == 38 && x == 17) || (y == 47 && x == 17) || (y == 15 && x == 18) || (y == 47 && x == 18) || (y == 47 && x == 19) || (y == 36 && x == 20) || (y == 37 && x == 20) || (y == 38 && x == 20) || (y == 39 && x == 20) || (y == 40 && x == 20) || (y == 41 && x == 20) || (y == 42 && x == 20) || (y == 43 && x == 20) || (y == 44 && x == 20) || (y == 45 && x == 20) || (y == 46 && x == 20) || (y == 47 && x == 20) || (y == 4 && x == 24) || (y == 5 && x == 24) || (y == 6 && x == 24) || (y == 7 && x == 24) || (y == 11 && x == 24) || (y == 12 && x == 24) || (y == 13 && x == 24) || (y == 14 && x == 24) || (y == 27 && x == 25) || (y == 27 && x == 26) || (y == 27 && x == 27) || (y == 41 && x == 27) || (y == 40 && x == 28) || (y == 21 && x == 29) || (y == 22 && x == 29) || (y == 30 && x == 29) || (y == 31 && x == 29) || (y == 37 && x == 31) || (y == 38 && x == 31) || (y == 39 && x == 31) || (y == 40 && x == 31) || (y == 41 && x == 31) || (y == 42 && x == 31) || (y == 43 && x == 31) || (y == 44 && x == 31) || (y == 45 && x == 31) || (y == 46 && x == 31) || (y == 47 && x == 31) || (y == 6 && x == 34) || (y == 7 && x == 34) || (y == 8 && x == 34) || (y == 9 && x == 34) || (y == 10 && x == 34) || (y == 11 && x == 34) || (y == 12 && x == 34) || (y == 13 && x == 34) || (y == 14 && x == 34) || (y == 39 && x == 36) || (y == 40 && x == 36) || (y == 44 && x == 36) || (y == 43 && x == 37)) oled_data <= 16'hb596;
        else if ((y == 41 && x == 14) || (y == 41 && x == 15)) oled_data <= 16'h18a2;
        else if ((y == 42 && x == 13) || (y == 10 && x == 20) || (y == 27 && x == 28)) oled_data <= 16'hef7d;
        else if ((y == 25 && x == 7) || (y == 25 && x == 17)) oled_data <= 16'h20e3;
        else if ((y == 46 && x == 10) || (y == 46 && x == 40)) oled_data <= 16'hb595;
        else if ((y == 12 && x == 27)) oled_data <= 16'h1021;
        else if ((y == 37 && x == 4) || (y == 5 && x == 30) || (y == 5 && x == 32) || (y == 37 && x == 34)) oled_data <= 16'h5a89;
        else if ((y == 8 && x == 24)) oled_data <= 16'had96;
        else if ((y == 25 && x == 19)) oled_data <= 16'h2061;
        else if ((y == 15 && x == 13) || (y == 9 && x == 15) || (y == 10 && x == 15) || (y == 40 && x == 25) || (y == 43 && x == 25) || (y == 44 && x == 25) || (y == 45 && x == 25) || (y == 46 && x == 25)) oled_data <= 16'hbdd7;
        else if ((y == 46 && x == 9) || (y == 46 && x == 39)) oled_data <= 16'h7bae;
        else if ((y == 26 && x == 17)) oled_data <= 16'hf7de;
        else if ((y == 39 && x == 9) || (y == 28 && x == 17) || (y == 39 && x == 39)) oled_data <= 16'h2903;
        else if ((y == 47 && x == 8) || (y == 47 && x == 38)) oled_data <= 16'h83cf;
        else if ((y == 41 && x == 9) || (y == 42 && x == 9) || (y == 41 && x == 39) || (y == 42 && x == 39)) oled_data <= 16'h3124;
        else if ((y == 23 && x == 18)) oled_data <= 16'h4a08;
        else if ((y == 20 && x == 22)) oled_data <= 16'ha513;
        else if ((y == 38 && x == 6) || (y == 6 && x == 30) || (y == 6 && x == 31) || (y == 38 && x == 36)) oled_data <= 16'h3186;
        else if ((y == 25 && x == 18)) oled_data <= 16'h49e7;
        else if ((y == 14 && x == 27)) oled_data <= 16'h6b4c;
        else if ((y == 47 && x == 4) || (y == 47 && x == 34)) oled_data <= 16'h49e8;
        else if ((y == 36 && x == 9) || (y == 36 && x == 39)) oled_data <= 16'h20e2;
        else if ((y == 5 && x == 15) || (y == 6 && x == 15) || (y == 8 && x == 15) || (y == 11 && x == 15) || (y == 13 && x == 15) || (y == 14 && x == 15) || (y == 47 && x == 29)) oled_data <= 16'had55;
        else if ((y == 27 && x == 17)) oled_data <= 16'h94b2;
        else if ((y == 6 && x == 6) || (y == 6 && x == 7) || (y == 6 && x == 8) || (y == 22 && x == 25) || (y == 37 && x == 25) || (y == 42 && x == 25) || (y == 22 && x == 26) || (y == 22 && x == 27) || (y == 22 && x == 28)) oled_data <= 16'hc618;
        else if ((y == 44 && x == 13) || (y == 30 && x == 23)) oled_data <= 16'hd699;
        else if ((y == 38 && x == 7) || (y == 38 && x == 37)) oled_data <= 16'h3986;
        else if ((y == 37 && x == 8) || (y == 4 && x == 28) || (y == 12 && x == 28) || (y == 13 && x == 28) || (y == 37 && x == 38)) oled_data <= 16'h8c30;
        else if ((y == 10 && x == 21)) oled_data <= 16'hce59;
        else if ((y == 25 && x == 8) || (y == 41 && x == 18) || (y == 41 && x == 19)) oled_data <= 16'h20a2;
        else if ((y == 37 && x == 9) || (y == 37 && x == 39)) oled_data <= 16'h6b4d;
        else if ((y == 10 && x == 22)) oled_data <= 16'hf73d;
        else if ((y == 37 && x == 6) || (y == 37 && x == 36)) oled_data <= 16'h5a8a;
        else if ((y == 7 && x == 15) || (y == 58 && x == 50)) oled_data <= 16'hb576;
        else if ((y == 42 && x == 15) || (y == 23 && x == 22) || (y == 24 && x == 22) || (y == 26 && x == 22) || (y == 27 && x == 22) || (y == 28 && x == 22) || (y == 29 && x == 22)) oled_data <= 16'ha4f3;
        else if ((y == 59 && x == 34)) oled_data <= 16'h7b6d;
        else if ((y == 38 && x == 8) || (y == 38 && x == 38)) oled_data <= 16'h73ae;
        else if ((y == 14 && x == 29)) oled_data <= 16'h6b2c;
        else if ((y == 10 && x == 18)) oled_data <= 16'hef5c;
        else if ((y == 38 && x == 5) || (y == 38 && x == 35)) oled_data <= 16'h3125;
        else if ((y == 39 && x == 8) || (y == 42 && x == 8) || (y == 45 && x == 8) || (y == 5 && x == 27) || (y == 39 && x == 38) || (y == 42 && x == 38) || (y == 45 && x == 38)) oled_data <= 16'h62eb;
        else if ((y == 31 && x == 23)) oled_data <= 16'hd6ba;
        else if ((y == 41 && x == 13)) oled_data <= 16'hd67a;
        else if ((y == 46 && x == 4) || (y == 46 && x == 5) || (y == 46 && x == 6) || (y == 46 && x == 7) || (y == 44 && x == 8) || (y == 14 && x == 30) || (y == 14 && x == 31) || (y == 14 && x == 32) || (y == 46 && x == 34) || (y == 46 && x == 35) || (y == 46 && x == 36) || (y == 46 && x == 37) || (y == 44 && x == 38) || (y == 59 && x == 43)) oled_data <= 16'h6aeb;
        else if ((y == 39 && x == 25)) oled_data <= 16'h83ee;
        else if ((y == 36 && x == 4) || (y == 36 && x == 6) || (y == 43 && x == 10) || (y == 21 && x == 19) || (y == 24 && x == 19) || (y == 4 && x == 30) || (y == 4 && x == 32) || (y == 36 && x == 34) || (y == 36 && x == 36) || (y == 43 && x == 40)) oled_data <= 16'h1820;
        else if ((y == 10 && x == 23) || (y == 23 && x == 23) || (y == 29 && x == 23) || (y == 42 && x == 30)) oled_data <= 16'hdeba;
        else if ((y == 23 && x == 6) || (y == 24 && x == 6) || (y == 29 && x == 6) || (y == 30 && x == 6)) oled_data <= 16'hce39;
        else if ((y == 43 && x == 8) || (y == 43 && x == 38)) oled_data <= 16'h732c;
        else if ((y == 22 && x == 11) || (y == 31 && x == 22) || (y == 55 && x == 41) || (y == 59 && x == 49) || (y == 55 && x == 56)) oled_data <= 16'hf7be;
        else if ((y == 26 && x == 16)) oled_data <= 16'hce58;
        else if ((y == 36 && x == 7) || (y == 36 && x == 37)) oled_data <= 16'h2021;
        else if ((y == 26 && x == 8) || (y == 42 && x == 18) || (y == 42 && x == 19) || (y == 25 && x == 22) || (y == 57 && x == 35) || (y == 57 && x == 48) || (y == 57 && x == 49)) oled_data <= 16'ha4d3;
        else if ((y == 15 && x == 27)) oled_data <= 16'h41e7;
        else if ((y == 20 && x == 17) || (y == 21 && x == 17) || (y == 22 && x == 17) || (y == 23 && x == 17) || (y == 29 && x == 17) || (y == 30 && x == 17) || (y == 55 && x == 45)) oled_data <= 16'h2924;
        else if ((y == 14 && x == 28)) oled_data <= 16'hb575;
        else if ((y == 6 && x == 4) || (y == 10 && x == 13) || (y == 26 && x == 13) || (y == 10 && x == 14) || (y == 26 && x == 19)) oled_data <= 16'hf77d;
        else if ((y == 5 && x == 33)) oled_data <= 16'h5aaa;
        else if ((y == 59 && x == 35)) oled_data <= 16'h8bf0;
        else if ((y == 5 && x == 4) || (y == 5 && x == 5) || (y == 5 && x == 6) || (y == 5 && x == 7) || (y == 27 && x == 7) || (y == 28 && x == 7) || (y == 5 && x == 8) || (y == 23 && x == 24) || (y == 21 && x == 25) || (y == 21 && x == 26) || (y == 8 && x == 27) || (y == 9 && x == 27) || (y == 10 && x == 27) || (y == 11 && x == 27) || (y == 21 && x == 27) || (y == 21 && x == 28) || (y == 12 && x == 29) || (y == 58 && x == 39) || (y == 58 && x == 45) || (y == 58 && x == 54)) oled_data <= 16'h1020;
        else if ((y == 38 && x == 9) || (y == 37 && x == 10) || (y == 38 && x == 39) || (y == 37 && x == 40)) oled_data <= 16'h5269;
        else if ((y == 44 && x == 9) || (y == 44 && x == 39)) oled_data <= 16'h3104;
        else if ((y == 4 && x == 4)) oled_data <= 16'h2040;
        else if ((y == 41 && x == 8) || (y == 47 && x == 9) || (y == 41 && x == 38) || (y == 47 && x == 39)) oled_data <= 16'h5acb;
        else if ((y == 36 && x == 31) || (y == 14 && x == 33)) oled_data <= 16'hb5b6;
        else if ((y == 15 && x == 28) || (y == 57 && x == 33) || (y == 57 && x == 34) || (y == 55 && x == 44)) oled_data <= 16'h9c92;
        else if ((y == 47 && x == 5) || (y == 47 && x == 6) || (y == 47 && x == 7) || (y == 15 && x == 29) || (y == 15 && x == 30) || (y == 15 && x == 31) || (y == 15 && x == 32) || (y == 47 && x == 35) || (y == 47 && x == 36) || (y == 47 && x == 37)) oled_data <= 16'h41e8;
        else if ((y == 26 && x == 6)) oled_data <= 16'heefc;
        else if ((y == 7 && x == 4) || (y == 7 && x == 28)) oled_data <= 16'h83ef;
        else if ((y == 21 && x == 22) || (y == 30 && x == 22)) oled_data <= 16'h9cf3;
        else if ((y == 10 && x == 19) || (y == 42 && x == 23) || (y == 22 && x == 24) || (y == 42 && x == 29)) oled_data <= 16'hef3c;
        else if ((y == 13 && x == 27) || (y == 54 && x == 44)) oled_data <= 16'h1040;
        else if ((y == 15 && x == 4) || (y == 15 && x == 5) || (y == 31 && x == 25) || (y == 31 && x == 26) || (y == 31 && x == 27) || (y == 31 && x == 28)) oled_data <= 16'hce79;
        else if ((y == 26 && x == 7) || (y == 42 && x == 14) || (y == 57 && x == 39) || (y == 57 && x == 54)) oled_data <= 16'h9cb2;
        else if ((y == 11 && x == 22) || (y == 38 && x == 25)) oled_data <= 16'h8bef;
        else if ((y == 23 && x == 7) || (y == 20 && x == 24)) oled_data <= 16'h820;
        else if ((y == 6 && x == 9) || (y == 26 && x == 15) || (y == 41 && x == 25)) oled_data <= 16'hc638;
        else if ((y == 26 && x == 18) || (y == 22 && x == 22)) oled_data <= 16'hef9d;
        else if ((y == 37 && x == 7) || (y == 5 && x == 31) || (y == 37 && x == 37)) oled_data <= 16'h5a69;
        else if ((y == 22 && x == 23)) oled_data <= 16'hffbe;
        else if ((y == 6 && x == 5) || (y == 25 && x == 28) || (y == 26 && x == 28)) oled_data <= 16'hef5d;
        else if ((y == 8 && x == 4) || (y == 9 && x == 4) || (y == 10 && x == 4) || (y == 11 && x == 4) || (y == 12 && x == 4) || (y == 13 && x == 4) || (y == 39 && x == 4) || (y == 9 && x == 5) || (y == 14 && x == 5) || (y == 20 && x == 5) || (y == 21 && x == 5) || (y == 41 && x == 5) || (y == 9 && x == 6) || (y == 9 && x == 7) || (y == 41 && x == 7) || (y == 42 && x == 7) || (y == 9 && x == 8) || (y == 24 && x == 8) || (y == 27 && x == 8) || (y == 5 && x == 9) || (y == 39 && x == 10) || (y == 40 && x == 10) || (y == 44 && x == 10) || (y == 45 && x == 10) || (y == 5 && x == 13) || (y == 8 && x == 13) || (y == 12 && x == 13) || (y == 21 && x == 13) || (y == 24 && x == 13) || (y == 28 && x == 13) || (y == 5 && x == 14) || (y == 8 && x == 14) || (y == 12 && x == 14) || (y == 21 && x == 14) || (y == 24 && x == 14) || (y == 28 && x == 14) || (y == 36 && x == 14) || (y == 37 && x == 14) || (y == 38 && x == 14) || (y == 39 && x == 14) || (y == 40 && x == 14) || (y == 44 && x == 14) || (y == 45 && x == 14) || (y == 46 && x == 14) || (y == 24 && x == 15) || (y == 36 && x == 15) || (y == 37 && x == 15) || (y == 38 && x == 15) || (y == 39 && x == 15) || (y == 40 && x == 15) || (y == 43 && x == 15) || (y == 44 && x == 15) || (y == 45 && x == 15) || (y == 46 && x == 15) || (y == 24 && x == 16) || (y == 7 && x == 18) || (y == 43 && x == 18) || (y == 4 && x == 19) || (y == 5 && x == 19) || (y == 8 && x == 19) || (y == 43 && x == 19) || (y == 12 && x == 20) || (y == 11 && x == 21) || (y == 7 && x == 22) || (y == 7 && x == 23) || (y == 8 && x == 23) || (y == 40 && x == 23) || (y == 43 && x == 23) || (y == 24 && x == 24) || (y == 25 && x == 24) || (y == 26 && x == 24) || (y == 27 && x == 24) || (y == 28 && x == 24) || (y == 29 && x == 24) || (y == 41 && x == 24) || (y == 44 && x == 24) || (y == 25 && x == 25) || (y == 30 && x == 25) || (y == 25 && x == 26) || (y == 26 && x == 26) || (y == 29 && x == 26) || (y == 30 && x == 26) || (y == 4 && x == 27) || (y == 25 && x == 27) || (y == 30 && x == 27) || (y == 39 && x == 27) || (y == 40 && x == 27) || (y == 30 && x == 28) || (y == 4 && x == 29) || (y == 7 && x == 29) || (y == 8 && x == 29) || (y == 9 && x == 29) || (y == 10 && x == 29) || (y == 11 && x == 29) || (y == 13 && x == 29) || (y == 40 && x == 29) || (y == 43 && x == 29) || (y == 39 && x == 30) || (y == 40 && x == 30) || (y == 7 && x == 32) || (y == 7 && x == 33) || (y == 59 && x == 33) || (y == 39 && x == 34) || (y == 41 && x == 35) || (y == 41 && x == 37) || (y == 42 && x == 37) || (y == 54 && x == 38) || (y == 39 && x == 40) || (y == 40 && x == 40) || (y == 44 && x == 40) || (y == 45 && x == 40) || (y == 57 && x == 44) || (y == 54 && x == 45) || (y == 56 && x == 45) || (y == 57 && x == 45) || (y == 54 && x == 53)) oled_data <= 16'h1000;
        else if ((y == 38 && x == 4) || (y == 6 && x == 32) || (y == 6 && x == 33) || (y == 38 && x == 34)) oled_data <= 16'h3145;
        else if ((y == 27 && x == 18) || (y == 5 && x == 28)) oled_data <= 16'ha514;
        else if ((y == 25 && x == 6)) oled_data <= 16'hc5f8;
        else if ((y == 5 && x == 29)) oled_data <= 16'h5268;
        else if ((y == 56 && x == 50)) oled_data <= 16'h2881;
        else if ((y == 59 && x == 45)) oled_data <= 16'h6b0b;
        else if ((y == 36 && x == 8) || (y == 36 && x == 38)) oled_data <= 16'h62aa;
        else if ((y == 40 && x == 8) || (y == 40 && x == 38)) oled_data <= 16'h62cb;
        else if ((y == 20 && x == 4) || (y == 21 && x == 4) || (y == 40 && x == 4) || (y == 41 && x == 4) || (y == 42 && x == 4) || (y == 43 && x == 4) || (y == 44 && x == 4) || (y == 45 && x == 4) || (y == 4 && x == 5) || (y == 10 && x == 5) || (y == 11 && x == 5) || (y == 12 && x == 5) || (y == 13 && x == 5) || (y == 36 && x == 5) || (y == 39 && x == 5) || (y == 40 && x == 5) || (y == 42 && x == 5) || (y == 43 && x == 5) || (y == 44 && x == 5) || (y == 45 && x == 5) || (y == 4 && x == 6) || (y == 10 && x == 6) || (y == 41 && x == 6) || (y == 42 && x == 6) || (y == 45 && x == 6) || (y == 4 && x == 7) || (y == 10 && x == 7) || (y == 45 && x == 7) || (y == 4 && x == 8) || (y == 10 && x == 8) || (y == 20 && x == 8) || (y == 21 && x == 8) || (y == 22 && x == 8) || (y == 23 && x == 8) || (y == 28 && x == 8) || (y == 29 && x == 8) || (y == 30 && x == 8) || (y == 4 && x == 9) || (y == 20 && x == 9) || (y == 21 && x == 9) || (y == 20 && x == 10) || (y == 21 && x == 10) || (y == 4 && x == 13) || (y == 6 && x == 13) || (y == 7 && x == 13) || (y == 9 && x == 13) || (y == 13 && x == 13) || (y == 14 && x == 13) || (y == 20 && x == 13) || (y == 22 && x == 13) || (y == 23 && x == 13) || (y == 25 && x == 13) || (y == 29 && x == 13) || (y == 30 && x == 13) || (y == 4 && x == 14) || (y == 6 && x == 14) || (y == 7 && x == 14) || (y == 9 && x == 14) || (y == 13 && x == 14) || (y == 14 && x == 14) || (y == 20 && x == 14) || (y == 22 && x == 14) || (y == 23 && x == 14) || (y == 25 && x == 14) || (y == 29 && x == 14) || (y == 30 && x == 14) || (y == 25 && x == 15) || (y == 36 && x == 16) || (y == 37 && x == 16) || (y == 45 && x == 16) || (y == 46 && x == 16) || (y == 36 && x == 17) || (y == 37 && x == 17) || (y == 45 && x == 17) || (y == 46 && x == 17) || (y == 4 && x == 18) || (y == 5 && x == 18) || (y == 6 && x == 18) || (y == 8 && x == 18) || (y == 12 && x == 18) || (y == 13 && x == 18) || (y == 14 && x == 18) || (y == 36 && x == 18) || (y == 37 && x == 18) || (y == 38 && x == 18) || (y == 39 && x == 18) || (y == 40 && x == 18) || (y == 44 && x == 18) || (y == 45 && x == 18) || (y == 46 && x == 18) || (y == 6 && x == 19) || (y == 7 && x == 19) || (y == 12 && x == 19) || (y == 13 && x == 19) || (y == 14 && x == 19) || (y == 20 && x == 19) || (y == 22 && x == 19) || (y == 23 && x == 19) || (y == 28 && x == 19) || (y == 29 && x == 19) || (y == 30 && x == 19) || (y == 36 && x == 19) || (y == 37 && x == 19) || (y == 38 && x == 19) || (y == 39 && x == 19) || (y == 40 && x == 19) || (y == 44 && x == 19) || (y == 45 && x == 19) || (y == 46 && x == 19) || (y == 12 && x == 21) || (y == 13 && x == 21) || (y == 4 && x == 22) || (y == 5 && x == 22) || (y == 6 && x == 22) || (y == 8 && x == 22) || (y == 12 && x == 22) || (y == 13 && x == 22) || (y == 14 && x == 22) || (y == 4 && x == 23) || (y == 5 && x == 23) || (y == 6 && x == 23) || (y == 11 && x == 23) || (y == 12 && x == 23) || (y == 13 && x == 23) || (y == 14 && x == 23) || (y == 36 && x == 23) || (y == 37 && x == 23) || (y == 38 && x == 23) || (y == 39 && x == 23) || (y == 41 && x == 23) || (y == 44 && x == 23) || (y == 45 && x == 23) || (y == 46 && x == 23) || (y == 37 && x == 24) || (y == 38 && x == 24) || (y == 40 && x == 24) || (y == 43 && x == 24) || (y == 45 && x == 24) || (y == 46 && x == 24) || (y == 20 && x == 25) || (y == 26 && x == 25) || (y == 29 && x == 25) || (y == 20 && x == 26) || (y == 20 && x == 27) || (y == 26 && x == 27) || (y == 29 && x == 27) || (y == 20 && x == 28) || (y == 29 && x == 28) || (y == 38 && x == 28) || (y == 39 && x == 28) || (y == 37 && x == 29) || (y == 38 && x == 29) || (y == 39 && x == 29) || (y == 41 && x == 29) || (y == 44 && x == 29) || (y == 45 && x == 29) || (y == 46 && x == 29) || (y == 13 && x == 30) || (y == 36 && x == 30) || (y == 37 && x == 30) || (y == 38 && x == 30) || (y == 43 && x == 30) || (y == 44 && x == 30) || (y == 45 && x == 30) || (y == 46 && x == 30) || (y == 4 && x == 31) || (y == 13 && x == 31) || (y == 8 && x == 32) || (y == 9 && x == 32) || (y == 10 && x == 32) || (y == 11 && x == 32) || (y == 12 && x == 32) || (y == 13 && x == 32) || (y == 8 && x == 33) || (y == 9 && x == 33) || (y == 10 && x == 33) || (y == 11 && x == 33) || (y == 12 && x == 33) || (y == 13 && x == 33) || (y == 54 && x == 33) || (y == 55 && x == 33) || (y == 56 && x == 33) || (y == 40 && x == 34) || (y == 41 && x == 34) || (y == 42 && x == 34) || (y == 43 && x == 34) || (y == 44 && x == 34) || (y == 45 && x == 34) || (y == 54 && x == 34) || (y == 56 && x == 34) || (y == 36 && x == 35) || (y == 39 && x == 35) || (y == 40 && x == 35) || (y == 42 && x == 35) || (y == 43 && x == 35) || (y == 44 && x == 35) || (y == 45 && x == 35) || (y == 54 && x == 35) || (y == 56 && x == 35) || (y == 58 && x == 35) || (y == 41 && x == 36) || (y == 42 && x == 36) || (y == 45 && x == 36) || (y == 45 && x == 37) || (y == 54 && x == 40) || (y == 56 && x == 43) || (y == 57 && x == 43) || (y == 58 && x == 43) || (y == 54 && x == 48) || (y == 55 && x == 48) || (y == 56 && x == 48) || (y == 58 && x == 48) || (y == 59 && x == 48) || (y == 54 && x == 49) || (y == 58 && x == 49) || (y == 54 && x == 50) || (y == 55 && x == 50) || (y == 59 && x == 50) || (y == 54 && x == 55)) oled_data <= 16'h1800;
        else if ((y == 36 && x == 13) || (y == 37 && x == 13) || (y == 38 && x == 13) || (y == 39 && x == 13) || (y == 40 && x == 13) || (y == 45 && x == 13) || (y == 46 && x == 13) || (y == 31 && x == 24)) oled_data <= 16'hd69a;
        else if ((y == 46 && x == 8) || (y == 46 && x == 38)) oled_data <= 16'h9cd2;
        else if ((y == 22 && x == 6)) oled_data <= 16'hbd96;
        else if (count <= 50_000_000) begin
            if ((y == 28 && x == 66) || (y == 44 && x == 66) || (y == 24 && x == 83) || (y == 27 && x == 85)) oled_data <= 16'h1062;
            else if ((y == 31 && x == 64) || (y == 41 && x == 64) || (y == 31 && x == 65) || (y == 32 && x == 68) || (y == 33 && x == 68) || (y == 34 && x == 68) || (y == 35 && x == 68) || (y == 36 && x == 68) || (y == 17 && x == 75) || (y == 18 && x == 75) || (y == 16 && x == 76) || (y == 16 && x == 77) || (y == 32 && x == 77) || (y == 33 && x == 77) || (y == 34 && x == 77) || (y == 35 && x == 77) || (y == 36 && x == 77) || (y == 16 && x == 78) || (y == 16 && x == 79) || (y == 16 && x == 80) || (y == 16 && x == 81)) oled_data <= 16'hef7d;
            else if ((y == 46 && x == 68) || (y == 47 && x == 79)) oled_data <= 16'h20e3;
            else if ((y == 30 && x == 70) || (y == 31 && x == 70) || (y == 30 && x == 71) || (y == 31 && x == 71) || (y == 32 && x == 71) || (y == 33 && x == 71) || (y == 34 && x == 71) || (y == 28 && x == 72) || (y == 29 && x == 72) || (y == 34 && x == 72) || (y == 35 && x == 72) || (y == 36 && x == 72) || (y == 28 && x == 73) || (y == 29 && x == 73) || (y == 34 && x == 73) || (y == 35 && x == 73) || (y == 36 && x == 73) || (y == 28 && x == 74) || (y == 29 && x == 74) || (y == 34 && x == 74) || (y == 35 && x == 74) || (y == 36 && x == 74) || (y == 28 && x == 75) || (y == 29 && x == 75) || (y == 34 && x == 75) || (y == 35 && x == 75) || (y == 36 && x == 75) || (y == 18 && x == 76) || (y == 19 && x == 76) || (y == 28 && x == 76) || (y == 29 && x == 76) || (y == 30 && x == 76) || (y == 31 && x == 76) || (y == 17 && x == 77) || (y == 18 && x == 77) || (y == 30 && x == 77) || (y == 31 && x == 77) || (y == 17 && x == 78) || (y == 20 && x == 78) || (y == 23 && x == 78) || (y == 30 && x == 78) || (y == 31 && x == 78) || (y == 32 && x == 78) || (y == 33 && x == 78) || (y == 34 && x == 78) || (y == 17 && x == 79) || (y == 23 && x == 79) || (y == 17 && x == 80) || (y == 18 && x == 80) || (y == 19 && x == 80) || (y == 23 && x == 80)) oled_data <= 16'h73af;
            else if ((y == 37 && x == 69) || (y == 37 && x == 76) || (y == 39 && x == 91) || (y == 39 && x == 92)) oled_data <= 16'hdeda;
            else if ((y == 35 && x == 71) || (y == 22 && x == 78) || (y == 35 && x == 78) || (y == 20 && x == 79) || (y == 22 && x == 79) || (y == 30 && x == 79) || (y == 31 && x == 79) || (y == 32 && x == 79) || (y == 33 && x == 79) || (y == 34 && x == 79) || (y == 22 && x == 80) || (y == 22 && x == 83)) oled_data <= 16'h630d;
            else if ((y == 22 && x == 72) || (y == 22 && x == 73) || (y == 20 && x == 76) || (y == 24 && x == 77) || (y == 24 && x == 78) || (y == 20 && x == 80) || (y == 22 && x == 84)) oled_data <= 16'h4a28;
            else if ((y == 48 && x == 81)) oled_data <= 16'h9c66;
            else if ((y == 47 && x == 67) || (y == 41 && x == 87) || (y == 42 && x == 87) || (y == 41 && x == 88) || (y == 42 && x == 88) || (y == 49 && x == 88) || (y == 44 && x == 90) || (y == 45 && x == 90) || (y == 46 && x == 90) || (y == 47 && x == 90)) oled_data <= 16'h3140;
            else if ((y == 52 && x == 81)) oled_data <= 16'hce57;
            else if ((y == 52 && x == 79) || (y == 37 && x == 93) || (y == 37 && x == 94)) oled_data <= 16'hb573;
            else if ((y == 45 && x == 80) || (y == 46 && x == 80) || (y == 30 && x == 91) || (y == 30 && x == 92)) oled_data <= 16'hb4a8;
            else if ((y == 39 && x == 68) || (y == 39 && x == 69) || (y == 35 && x == 70) || (y == 37 && x == 72) || (y == 37 && x == 73) || (y == 37 && x == 74) || (y == 37 && x == 75) || (y == 24 && x == 76) || (y == 39 && x == 76) || (y == 20 && x == 77) || (y == 39 && x == 77) || (y == 35 && x == 79) || (y == 23 && x == 83)) oled_data <= 16'h528a;
            else if ((y == 49 && x == 69) || (y == 50 && x == 77) || (y == 49 && x == 78) || (y == 47 && x == 81) || (y == 42 && x == 82) || (y == 43 && x == 82) || (y == 44 && x == 82) || (y == 49 && x == 82) || (y == 31 && x == 92) || (y == 32 && x == 93) || (y == 32 && x == 94)) oled_data <= 16'hb4a6;
            else if ((y == 29 && x == 66) || (y == 30 && x == 66) || (y == 31 && x == 66) || (y == 41 && x == 66) || (y == 42 && x == 66) || (y == 43 && x == 66) || (y == 27 && x == 68) || (y == 45 && x == 68) || (y == 24 && x == 70) || (y == 46 && x == 72)) oled_data <= 16'h2104;
            else if ((y == 47 && x == 66) || (y == 50 && x == 88) || (y == 48 && x == 90)) oled_data <= 16'h4a04;
            else if ((y == 37 && x == 67) || (y == 38 && x == 67) || (y == 30 && x == 68) || (y == 40 && x == 68) || (y == 30 && x == 69) || (y == 31 && x == 69) || (y == 40 && x == 69) || (y == 28 && x == 70) || (y == 29 && x == 70) || (y == 39 && x == 70) || (y == 40 && x == 70) || (y == 41 && x == 70) || (y == 42 && x == 70) || (y == 24 && x == 71) || (y == 28 && x == 71) || (y == 36 && x == 71) || (y == 37 && x == 71) || (y == 38 && x == 71) || (y == 39 && x == 71) || (y == 40 && x == 71) || (y == 41 && x == 71) || (y == 42 && x == 71) || (y == 26 && x == 72) || (y == 27 && x == 72) || (y == 38 && x == 72) || (y == 39 && x == 72) || (y == 40 && x == 72) || (y == 41 && x == 72) || (y == 42 && x == 72) || (y == 43 && x == 72) || (y == 44 && x == 72) || (y == 26 && x == 73) || (y == 27 && x == 73) || (y == 38 && x == 73) || (y == 39 && x == 73) || (y == 40 && x == 73) || (y == 41 && x == 73) || (y == 42 && x == 73) || (y == 43 && x == 73) || (y == 44 && x == 73) || (y == 24 && x == 74) || (y == 26 && x == 74) || (y == 27 && x == 74) || (y == 38 && x == 74) || (y == 39 && x == 74) || (y == 40 && x == 74) || (y == 41 && x == 74) || (y == 42 && x == 74) || (y == 43 && x == 74) || (y == 44 && x == 74) || (y == 24 && x == 75) || (y == 26 && x == 75) || (y == 27 && x == 75) || (y == 38 && x == 75) || (y == 39 && x == 75) || (y == 40 && x == 75) || (y == 41 && x == 75) || (y == 42 && x == 75) || (y == 43 && x == 75) || (y == 44 && x == 75) || (y == 25 && x == 76) || (y == 26 && x == 76) || (y == 27 && x == 76) || (y == 40 && x == 76) || (y == 41 && x == 76) || (y == 42 && x == 76) || (y == 43 && x == 76) || (y == 44 && x == 76) || (y == 25 && x == 77) || (y == 26 && x == 77) || (y == 27 && x == 77) || (y == 40 && x == 77) || (y == 41 && x == 77) || (y == 42 && x == 77) || (y == 43 && x == 77) || (y == 44 && x == 77) || (y == 25 && x == 78) || (y == 26 && x == 78) || (y == 27 && x == 78) || (y == 28 && x == 78) || (y == 29 && x == 78) || (y == 36 && x == 78) || (y == 37 && x == 78) || (y == 38 && x == 78) || (y == 39 && x == 78) || (y == 40 && x == 78) || (y == 41 && x == 78) || (y == 42 && x == 78) || (y == 43 && x == 78) || (y == 44 && x == 78) || (y == 24 && x == 79) || (y == 26 && x == 79) || (y == 27 && x == 79) || (y == 28 && x == 79) || (y == 29 && x == 79) || (y == 36 && x == 79) || (y == 37 && x == 79) || (y == 38 && x == 79) || (y == 39 && x == 79) || (y == 40 && x == 79) || (y == 41 && x == 79) || (y == 42 && x == 79) || (y == 26 && x == 80) || (y == 27 && x == 80) || (y == 28 && x == 80) || (y == 29 && x == 80) || (y == 30 && x == 80) || (y == 31 && x == 80) || (y == 32 && x == 80) || (y == 33 && x == 80) || (y == 34 && x == 80) || (y == 35 && x == 80) || (y == 36 && x == 80) || (y == 37 && x == 80) || (y == 38 && x == 80) || (y == 39 && x == 80) || (y == 40 && x == 80) || (y == 41 && x == 80) || (y == 42 && x == 80) || (y == 28 && x == 81) || (y == 29 && x == 81) || (y == 30 && x == 81) || (y == 31 && x == 81) || (y == 32 && x == 81) || (y == 33 && x == 81) || (y == 34 && x == 81) || (y == 35 && x == 81) || (y == 36 && x == 81) || (y == 37 && x == 81) || (y == 38 && x == 81) || (y == 39 && x == 81) || (y == 40 && x == 81) || (y == 24 && x == 82) || (y == 28 && x == 82) || (y == 29 && x == 82) || (y == 30 && x == 82) || (y == 31 && x == 82) || (y == 32 && x == 82) || (y == 33 && x == 82) || (y == 34 && x == 82) || (y == 35 && x == 82) || (y == 36 && x == 82) || (y == 37 && x == 82) || (y == 38 && x == 82) || (y == 39 && x == 82) || (y == 40 && x == 82) || (y == 28 && x == 83) || (y == 29 && x == 83) || (y == 30 && x == 83) || (y == 31 && x == 83) || (y == 32 && x == 83) || (y == 33 && x == 83) || (y == 34 && x == 83) || (y == 35 && x == 83) || (y == 36 && x == 83) || (y == 37 && x == 83) || (y == 38 && x == 83) || (y == 28 && x == 84) || (y == 29 && x == 84) || (y == 30 && x == 84) || (y == 31 && x == 84) || (y == 32 && x == 84) || (y == 33 && x == 84) || (y == 34 && x == 84) || (y == 35 && x == 84) || (y == 36 && x == 84) || (y == 37 && x == 84) || (y == 38 && x == 84) || (y == 32 && x == 85) || (y == 33 && x == 85) || (y == 34 && x == 85) || (y == 35 && x == 85) || (y == 36 && x == 85) || (y == 32 && x == 86) || (y == 33 && x == 86) || (y == 34 && x == 86) || (y == 35 && x == 86) || (y == 36 && x == 86)) oled_data <= 16'h39a7;
            else if ((y == 49 && x == 87) || (y == 44 && x == 89) || (y == 45 && x == 89) || (y == 46 && x == 89) || (y == 47 && x == 89)) oled_data <= 16'h3940;
            else if ((y == 50 && x == 79) || (y == 49 && x == 81) || (y == 50 && x == 81)) oled_data <= 16'h8b86;
            else if ((y == 33 && x == 65) || (y == 34 && x == 65) || (y == 35 && x == 65) || (y == 36 && x == 65) || (y == 37 && x == 65) || (y == 38 && x == 65) || (y == 39 && x == 65) || (y == 29 && x == 67) || (y == 30 && x == 67) || (y == 31 && x == 67) || (y == 41 && x == 67) || (y == 42 && x == 67) || (y == 43 && x == 67) || (y == 26 && x == 68) || (y == 27 && x == 69) || (y == 45 && x == 69) || (y == 45 && x == 70) || (y == 25 && x == 71) || (y == 45 && x == 71) || (y == 25 && x == 72) || (y == 25 && x == 73) || (y == 47 && x == 73) || (y == 47 && x == 74) || (y == 21 && x == 75) || (y == 47 && x == 75) || (y == 21 && x == 76) || (y == 47 && x == 76) || (y == 21 && x == 77) || (y == 47 && x == 77) || (y == 21 && x == 78) || (y == 47 && x == 78) || (y == 21 && x == 79) || (y == 21 && x == 80) || (y == 21 && x == 81) || (y == 21 && x == 82) || (y == 25 && x == 82) || (y == 25 && x == 83) || (y == 29 && x == 87) || (y == 30 && x == 87) || (y == 31 && x == 87) || (y == 39 && x == 87) || (y == 30 && x == 88) || (y == 31 && x == 88) || (y == 31 && x == 89) || (y == 32 && x == 89) || (y == 33 && x == 89) || (y == 34 && x == 89) || (y == 35 && x == 89) || (y == 36 && x == 89) || (y == 37 && x == 89) || (y == 38 && x == 89) || (y == 38 && x == 90)) oled_data <= 16'h841;
            else if ((y == 48 && x == 73) || (y == 48 && x == 79) || (y == 43 && x == 89) || (y == 34 && x == 94) || (y == 35 && x == 94) || (y == 36 && x == 94)) oled_data <= 16'h2900;
            else if ((y == 49 && x == 74) || (y == 49 && x == 75) || (y == 49 && x == 76) || (y == 49 && x == 85) || (y == 49 && x == 86) || (y == 45 && x == 87) || (y == 46 && x == 87) || (y == 47 && x == 87) || (y == 45 && x == 88) || (y == 46 && x == 88)) oled_data <= 16'hdd85;
            else if ((y == 47 && x == 68) || (y == 42 && x == 83) || (y == 43 && x == 83) || (y == 44 && x == 83) || (y == 49 && x == 83) || (y == 41 && x == 84) || (y == 41 && x == 85) || (y == 41 && x == 86) || (y == 33 && x == 92)) oled_data <= 16'hee88;
            else if ((y == 32 && x == 66) || (y == 33 && x == 66) || (y == 39 && x == 66) || (y == 40 && x == 66) || (y == 32 && x == 67) || (y == 33 && x == 67) || (y == 40 && x == 67) || (y == 28 && x == 68) || (y == 41 && x == 68) || (y == 42 && x == 68) || (y == 43 && x == 68) || (y == 44 && x == 68) || (y == 28 && x == 69) || (y == 29 && x == 69) || (y == 42 && x == 69) || (y == 43 && x == 69) || (y == 44 && x == 69) || (y == 26 && x == 70) || (y == 27 && x == 70) || (y == 43 && x == 70) || (y == 44 && x == 70) || (y == 26 && x == 71) || (y == 27 && x == 71) || (y == 43 && x == 71) || (y == 44 && x == 71) || (y == 45 && x == 72) || (y == 45 && x == 73) || (y == 46 && x == 73) || (y == 25 && x == 74) || (y == 45 && x == 74) || (y == 46 && x == 74) || (y == 25 && x == 75) || (y == 45 && x == 75) || (y == 46 && x == 75) || (y == 45 && x == 76) || (y == 46 && x == 76) || (y == 45 && x == 77) || (y == 46 && x == 77) || (y == 45 && x == 78) || (y == 46 && x == 78) || (y == 25 && x == 80) || (y == 43 && x == 80) || (y == 26 && x == 82) || (y == 27 && x == 82) || (y == 26 && x == 83) || (y == 27 && x == 83) || (y == 26 && x == 84) || (y == 27 && x == 84) || (y == 28 && x == 86) || (y == 29 && x == 86) || (y == 30 && x == 86) || (y == 31 && x == 86) || (y == 38 && x == 86) || (y == 32 && x == 87) || (y == 33 && x == 87) || (y == 34 && x == 87) || (y == 35 && x == 87) || (y == 36 && x == 87) || (y == 37 && x == 87) || (y == 38 && x == 87) || (y == 32 && x == 88) || (y == 33 && x == 88) || (y == 34 && x == 88) || (y == 35 && x == 88) || (y == 36 && x == 88) || (y == 37 && x == 88) || (y == 38 && x == 88)) oled_data <= 16'h20e5;
            else if ((y == 48 && x == 68) || (y == 50 && x == 70) || (y == 50 && x == 71) || (y == 50 && x == 72) || (y == 50 && x == 73) || (y == 46 && x == 81) || (y == 50 && x == 84)) oled_data <= 16'hde26;
            else if ((y == 49 && x == 77) || (y == 47 && x == 88) || (y == 34 && x == 91) || (y == 35 && x == 91) || (y == 36 && x == 91) || (y == 34 && x == 92) || (y == 35 && x == 92) || (y == 36 && x == 92)) oled_data <= 16'hdd87;
            else if ((y == 39 && x == 83)) oled_data <= 16'h39a5;
            else if ((y == 32 && x == 70) || (y == 33 && x == 70) || (y == 34 && x == 70) || (y == 17 && x == 76) || (y == 28 && x == 77) || (y == 29 && x == 77) || (y == 20 && x == 81)) oled_data <= 16'h6b6e;
            else if ((y == 48 && x == 72) || (y == 48 && x == 74) || (y == 48 && x == 75) || (y == 48 && x == 76) || (y == 48 && x == 77) || (y == 48 && x == 78) || (y == 43 && x == 90)) oled_data <= 16'h20a0;
            else if ((y == 30 && x == 72) || (y == 31 && x == 72) || (y == 32 && x == 72) || (y == 33 && x == 72) || (y == 30 && x == 73) || (y == 31 && x == 73) || (y == 32 && x == 73) || (y == 33 && x == 73) || (y == 23 && x == 74) || (y == 30 && x == 74) || (y == 31 && x == 74) || (y == 32 && x == 74) || (y == 33 && x == 74) || (y == 23 && x == 75) || (y == 30 && x == 75) || (y == 31 && x == 75) || (y == 32 && x == 75) || (y == 33 && x == 75) || (y == 22 && x == 76)) oled_data <= 16'h94f3;
            else if ((y == 32 && x == 65) || (y == 40 && x == 65) || (y == 28 && x == 67) || (y == 44 && x == 67) || (y == 26 && x == 69) || (y == 46 && x == 69) || (y == 25 && x == 70) || (y == 46 && x == 70) || (y == 46 && x == 71) || (y == 23 && x == 72) || (y == 47 && x == 72) || (y == 23 && x == 73) || (y == 21 && x == 74) || (y == 26 && x == 85) || (y == 26 && x == 86) || (y == 28 && x == 87) || (y == 40 && x == 87) || (y == 28 && x == 88) || (y == 29 && x == 88) || (y == 39 && x == 88) || (y == 40 && x == 88) || (y == 30 && x == 89) || (y == 30 && x == 90) || (y == 31 && x == 90) || (y == 32 && x == 90) || (y == 33 && x == 90) || (y == 34 && x == 90) || (y == 35 && x == 90) || (y == 36 && x == 90) || (y == 37 && x == 90)) oled_data <= 16'h0;
            else if ((y == 50 && x == 74) || (y == 50 && x == 75) || (y == 50 && x == 76) || (y == 50 && x == 85) || (y == 50 && x == 86) || (y == 48 && x == 87) || (y == 48 && x == 88) || (y == 31 && x == 91)) oled_data <= 16'hc4e6;
            else if ((y == 50 && x == 66) || (y == 51 && x == 79)) oled_data <= 16'h6b0a;
            else if ((y == 48 && x == 67) || (y == 49 && x == 67) || (y == 51 && x == 69) || (y == 51 && x == 70) || (y == 51 && x == 71) || (y == 51 && x == 72) || (y == 51 && x == 73) || (y == 51 && x == 74) || (y == 51 && x == 75) || (y == 51 && x == 76) || (y == 51 && x == 77) || (y == 51 && x == 78) || (y == 47 && x == 80) || (y == 48 && x == 80) || (y == 49 && x == 80) || (y == 51 && x == 82) || (y == 51 && x == 83) || (y == 40 && x == 84) || (y == 51 && x == 84) || (y == 40 && x == 85) || (y == 51 && x == 85) || (y == 40 && x == 86) || (y == 51 && x == 86) || (y == 38 && x == 91) || (y == 38 && x == 92) || (y == 34 && x == 93) || (y == 35 && x == 93) || (y == 36 && x == 93)) oled_data <= 16'h39a2;
            else if ((y == 52 && x == 68) || (y == 52 && x == 69) || (y == 52 && x == 70) || (y == 52 && x == 71) || (y == 52 && x == 72) || (y == 52 && x == 73) || (y == 52 && x == 74) || (y == 52 && x == 75) || (y == 52 && x == 76) || (y == 52 && x == 77) || (y == 52 && x == 78) || (y == 51 && x == 81) || (y == 52 && x == 82) || (y == 52 && x == 83) || (y == 52 && x == 84) || (y == 52 && x == 85) || (y == 52 && x == 86)) oled_data <= 16'h9490;
            else if ((y == 48 && x == 69) || (y == 45 && x == 82) || (y == 48 && x == 82) || (y == 48 && x == 83) || (y == 48 && x == 85) || (y == 48 && x == 86) || (y == 43 && x == 87) || (y == 32 && x == 91) || (y == 33 && x == 91) || (y == 32 && x == 92)) oled_data <= 16'hfec6;
            else if ((y == 48 && x == 66) || (y == 49 && x == 66) || (y == 50 && x == 67) || (y == 51 && x == 68) || (y == 45 && x == 79) || (y == 46 && x == 79) || (y == 50 && x == 80)) oled_data <= 16'h5246;
            else if ((y == 37 && x == 91) || (y == 37 && x == 92)) oled_data <= 16'h8363;
            else if ((y == 40 && x == 83) || (y == 39 && x == 84) || (y == 39 && x == 85) || (y == 39 && x == 86)) oled_data <= 16'h39a4;
            else if ((y == 34 && x == 66) || (y == 35 && x == 66) || (y == 36 && x == 66) || (y == 37 && x == 66) || (y == 38 && x == 66) || (y == 34 && x == 67) || (y == 35 && x == 67) || (y == 36 && x == 67) || (y == 31 && x == 68) || (y == 29 && x == 71) || (y == 25 && x == 79) || (y == 43 && x == 79) || (y == 44 && x == 79) || (y == 24 && x == 81)) oled_data <= 16'h3166;
            else if ((y == 47 && x == 69) || (y == 47 && x == 70) || (y == 48 && x == 70) || (y == 49 && x == 70) || (y == 47 && x == 71) || (y == 48 && x == 71) || (y == 49 && x == 71) || (y == 49 && x == 72) || (y == 49 && x == 73) || (y == 46 && x == 82) || (y == 47 && x == 82) || (y == 45 && x == 83) || (y == 46 && x == 83) || (y == 47 && x == 83) || (y == 42 && x == 84) || (y == 43 && x == 84) || (y == 44 && x == 84) || (y == 45 && x == 84) || (y == 46 && x == 84) || (y == 47 && x == 84) || (y == 48 && x == 84) || (y == 49 && x == 84) || (y == 42 && x == 85) || (y == 43 && x == 85) || (y == 44 && x == 85) || (y == 45 && x == 85) || (y == 46 && x == 85) || (y == 47 && x == 85) || (y == 42 && x == 86) || (y == 43 && x == 86) || (y == 44 && x == 86) || (y == 45 && x == 86) || (y == 46 && x == 86) || (y == 47 && x == 86) || (y == 44 && x == 87) || (y == 44 && x == 88)) oled_data <= 16'hff05;
            else if ((y == 43 && x == 88)) oled_data <= 16'hff2a;
            else if ((y == 31 && x == 93) || (y == 31 && x == 94)) oled_data <= 16'hef39;
            else if ((y == 37 && x == 70) || (y == 38 && x == 70) || (y == 24 && x == 80) || (y == 26 && x == 81) || (y == 27 && x == 81) || (y == 37 && x == 85) || (y == 37 && x == 86)) oled_data <= 16'h3146;
            else if ((y == 29 && x == 68) || (y == 44 && x == 80) || (y == 25 && x == 81)) oled_data <= 16'h18c4;
            else if ((y == 24 && x == 72) || (y == 24 && x == 73) || (y == 23 && x == 84) || (y == 24 && x == 84) || (y == 25 && x == 84) || (y == 27 && x == 86)) oled_data <= 16'h800;
            else if ((y == 50 && x == 64) || (y == 46 && x == 66) || (y == 51 && x == 87) || (y == 52 && x == 87) || (y == 41 && x == 89) || (y == 42 && x == 89) || (y == 49 && x == 89) || (y == 50 && x == 89) || (y == 29 && x == 91) || (y == 29 && x == 92)) oled_data <= 16'hffde;
            else if ((y == 32 && x == 64) || (y == 33 && x == 64) || (y == 34 && x == 64) || (y == 35 && x == 64) || (y == 36 && x == 64) || (y == 37 && x == 64) || (y == 38 && x == 64) || (y == 39 && x == 64) || (y == 40 && x == 64) || (y == 22 && x == 74) || (y == 22 && x == 75) || (y == 19 && x == 77) || (y == 18 && x == 79)) oled_data <= 16'h7bef;
            else if ((y == 41 && x == 81)) oled_data <= 16'h83aa;
            else if ((y == 50 && x == 87) || (y == 48 && x == 89)) oled_data <= 16'h5a64;
            else if ((y == 49 && x == 68) || (y == 50 && x == 68) || (y == 50 && x == 69) || (y == 50 && x == 78) || (y == 49 && x == 79) || (y == 41 && x == 82) || (y == 50 && x == 82) || (y == 33 && x == 93) || (y == 33 && x == 94)) oled_data <= 16'ha447;
            else if ((y == 38 && x == 69) || (y == 23 && x == 76) || (y == 38 && x == 76) || (y == 23 && x == 77) || (y == 37 && x == 77) || (y == 19 && x == 78) || (y == 23 && x == 81) || (y == 22 && x == 82) || (y == 21 && x == 83)) oled_data <= 16'hce59;
            else if ((y == 42 && x == 81) || (y == 43 && x == 81) || (y == 44 && x == 81)) oled_data <= 16'h7305;
            else if ((y == 41 && x == 65) || (y == 37 && x == 68) || (y == 20 && x == 83) || (y == 22 && x == 85) || (y == 23 && x == 85) || (y == 24 && x == 85) || (y == 25 && x == 85) || (y == 39 && x == 89) || (y == 39 && x == 90)) oled_data <= 16'hd69a;
            else if ((y == 39 && x == 67) || (y == 41 && x == 69) || (y == 36 && x == 70) || (y == 28 && x == 85) || (y == 29 && x == 85) || (y == 30 && x == 85) || (y == 31 && x == 85) || (y == 38 && x == 85)) oled_data <= 16'h2905;
            else if ((y == 20 && x == 74) || (y == 20 && x == 75) || (y == 22 && x == 77) || (y == 18 && x == 78) || (y == 22 && x == 81) || (y == 20 && x == 82)) oled_data <= 16'h8c92;
            else if ((y == 38 && x == 68) || (y == 38 && x == 77) || (y == 19 && x == 79) || (y == 17 && x == 81) || (y == 18 && x == 81) || (y == 19 && x == 81)) oled_data <= 16'hb5b6;
            else if ((y == 45 && x == 81) || (y == 41 && x == 83) || (y == 50 && x == 83)) oled_data <= 16'hd5e8;
            else oled_data <= 16'hffff; 
        end
        else if (count <= 100_000_000) begin
            if ((y == 17 && x == 81)) oled_data <= 16'hf529;
            else if ((y == 27 && x == 66) || (y == 43 && x == 66) || (y == 23 && x == 83) || (y == 26 && x == 85) || (y == 38 && x == 87)) oled_data <= 16'h1062;
            else if ((y == 36 && x == 69) || (y == 36 && x == 76) || (y == 38 && x == 91) || (y == 38 && x == 92)) oled_data <= 16'hdeda;
            else if ((y == 21 && x == 72) || (y == 21 && x == 73) || (y == 23 && x == 77) || (y == 21 && x == 84)) oled_data <= 16'h4a28;
            else if ((y == 46 && x == 67) || (y == 44 && x == 87) || (y == 45 && x == 88) || (y == 46 && x == 88) || (y == 47 && x == 88) || (y == 48 && x == 88)) oled_data <= 16'h3140;
            else if ((y == 42 && x == 82) || (y == 42 && x == 83) || (y == 42 && x == 84) || (y == 29 && x == 91) || (y == 29 && x == 92)) oled_data <= 16'hb4a8;
            else if ((y == 38 && x == 68) || (y == 38 && x == 69) || (y == 34 && x == 70) || (y == 36 && x == 72) || (y == 36 && x == 73) || (y == 36 && x == 74) || (y == 36 && x == 75) || (y == 23 && x == 76) || (y == 38 && x == 76) || (y == 38 && x == 77) || (y == 34 && x == 79)) oled_data <= 16'h528a;
            else if ((y == 17 && x == 82)) oled_data <= 16'hf50c;
            else if ((y == 32 && x == 65) || (y == 33 && x == 65) || (y == 34 && x == 65) || (y == 35 && x == 65) || (y == 36 && x == 65) || (y == 37 && x == 65) || (y == 38 && x == 65) || (y == 28 && x == 67) || (y == 29 && x == 67) || (y == 30 && x == 67) || (y == 40 && x == 67) || (y == 41 && x == 67) || (y == 42 && x == 67) || (y == 25 && x == 68) || (y == 26 && x == 69) || (y == 44 && x == 69) || (y == 44 && x == 70) || (y == 24 && x == 71) || (y == 44 && x == 71) || (y == 24 && x == 72) || (y == 24 && x == 73) || (y == 46 && x == 73) || (y == 20 && x == 75) || (y == 20 && x == 76) || (y == 20 && x == 77) || (y == 20 && x == 78) || (y == 20 && x == 79) || (y == 20 && x == 80) || (y == 20 && x == 81) || (y == 20 && x == 82) || (y == 24 && x == 82) || (y == 24 && x == 83) || (y == 28 && x == 87) || (y == 29 && x == 87) || (y == 30 && x == 87) || (y == 39 && x == 87) || (y == 40 && x == 87) || (y == 29 && x == 88) || (y == 30 && x == 88) || (y == 30 && x == 89) || (y == 31 && x == 89) || (y == 32 && x == 89) || (y == 33 && x == 89) || (y == 34 && x == 89) || (y == 35 && x == 89) || (y == 36 && x == 89) || (y == 37 && x == 89) || (y == 37 && x == 90)) oled_data <= 16'h841;
            else if ((y == 48 && x == 78) || (y == 48 && x == 84) || (y == 46 && x == 85) || (y == 47 && x == 85)) oled_data <= 16'hdd85;
            else if ((y == 42 && x == 77) || (y == 43 && x == 77)) oled_data <= 16'h39a5;
            else if ((y == 31 && x == 65) || (y == 39 && x == 65) || (y == 27 && x == 67) || (y == 43 && x == 67) || (y == 25 && x == 69) || (y == 45 && x == 69) || (y == 24 && x == 70) || (y == 45 && x == 70) || (y == 45 && x == 71) || (y == 22 && x == 72) || (y == 46 && x == 72) || (y == 22 && x == 73) || (y == 20 && x == 74) || (y == 24 && x == 84) || (y == 25 && x == 85) || (y == 25 && x == 86) || (y == 27 && x == 87) || (y == 41 && x == 87) || (y == 27 && x == 88) || (y == 28 && x == 88) || (y == 38 && x == 88) || (y == 39 && x == 88) || (y == 40 && x == 88) || (y == 41 && x == 88) || (y == 29 && x == 89) || (y == 29 && x == 90) || (y == 30 && x == 90) || (y == 31 && x == 90) || (y == 32 && x == 90) || (y == 33 && x == 90) || (y == 34 && x == 90) || (y == 35 && x == 90) || (y == 36 && x == 90)) oled_data <= 16'h0;
            else if ((y == 48 && x == 77) || (y == 49 && x == 78) || (y == 49 && x == 84) || (y == 48 && x == 85) || (y == 30 && x == 91)) oled_data <= 16'hc4e6;
            else if ((y == 51 && x == 68) || (y == 51 && x == 69) || (y == 51 && x == 70) || (y == 51 && x == 71) || (y == 51 && x == 72) || (y == 51 && x == 73) || (y == 51 && x == 74) || (y == 51 && x == 75) || (y == 51 && x == 76) || (y == 51 && x == 77) || (y == 51 && x == 78) || (y == 51 && x == 79) || (y == 51 && x == 80) || (y == 51 && x == 81) || (y == 51 && x == 82) || (y == 51 && x == 83) || (y == 51 && x == 84) || (y == 51 && x == 85) || (y == 51 && x == 86)) oled_data <= 16'h9490;
            else if ((y == 15 && x == 83)) oled_data <= 16'hec85;
            else if ((y == 24 && x == 81)) oled_data <= 16'h18c4;
            else if ((y == 23 && x == 72) || (y == 23 && x == 73) || (y == 22 && x == 84) || (y == 23 && x == 84) || (y == 26 && x == 86)) oled_data <= 16'h800;
            else if ((y == 45 && x == 66) || (y == 15 && x == 75) || (y == 13 && x == 77) || (y == 11 && x == 80) || (y == 11 && x == 81) || (y == 11 && x == 82) || (y == 13 && x == 85) || (y == 42 && x == 87) || (y == 50 && x == 87) || (y == 51 && x == 87) || (y == 44 && x == 89) || (y == 45 && x == 89) || (y == 46 && x == 89) || (y == 47 && x == 89) || (y == 48 && x == 89) || (y == 49 && x == 89) || (y == 28 && x == 91) || (y == 28 && x == 92)) oled_data <= 16'hffde;
            else if ((y == 42 && x == 85) || (y == 49 && x == 87)) oled_data <= 16'h5a64;
            else if ((y == 48 && x == 68) || (y == 49 && x == 68) || (y == 49 && x == 69) || (y == 49 && x == 76) || (y == 49 && x == 86) || (y == 32 && x == 93) || (y == 32 && x == 94)) oled_data <= 16'ha447;
            else if ((y == 13 && x == 78) || (y == 13 && x == 84)) oled_data <= 16'hffbd;
            else if ((y == 40 && x == 64) || (y == 30 && x == 65) || (y == 31 && x == 68) || (y == 32 && x == 68) || (y == 33 && x == 68) || (y == 34 && x == 68) || (y == 35 && x == 68) || (y == 31 && x == 77) || (y == 32 && x == 77) || (y == 33 && x == 77) || (y == 34 && x == 77) || (y == 35 && x == 77)) oled_data <= 16'hef7d;
            else if ((y == 45 && x == 68) || (y == 45 && x == 75)) oled_data <= 16'h20e3;
            else if ((y == 29 && x == 70) || (y == 30 && x == 70) || (y == 29 && x == 71) || (y == 30 && x == 71) || (y == 31 && x == 71) || (y == 32 && x == 71) || (y == 33 && x == 71) || (y == 27 && x == 72) || (y == 28 && x == 72) || (y == 33 && x == 72) || (y == 34 && x == 72) || (y == 35 && x == 72) || (y == 27 && x == 73) || (y == 28 && x == 73) || (y == 33 && x == 73) || (y == 34 && x == 73) || (y == 35 && x == 73) || (y == 27 && x == 74) || (y == 28 && x == 74) || (y == 33 && x == 74) || (y == 34 && x == 74) || (y == 35 && x == 74) || (y == 27 && x == 75) || (y == 28 && x == 75) || (y == 33 && x == 75) || (y == 34 && x == 75) || (y == 35 && x == 75) || (y == 27 && x == 76) || (y == 28 && x == 76) || (y == 29 && x == 76) || (y == 30 && x == 76) || (y == 29 && x == 77) || (y == 30 && x == 77) || (y == 22 && x == 78) || (y == 29 && x == 78) || (y == 30 && x == 78) || (y == 31 && x == 78) || (y == 32 && x == 78) || (y == 33 && x == 78) || (y == 22 && x == 79) || (y == 22 && x == 80)) oled_data <= 16'h73af;
            else if ((y == 28 && x == 66) || (y == 29 && x == 66) || (y == 30 && x == 66) || (y == 40 && x == 66) || (y == 41 && x == 66) || (y == 42 && x == 66) || (y == 26 && x == 68) || (y == 44 && x == 68) || (y == 23 && x == 70) || (y == 45 && x == 72) || (y == 45 && x == 74) || (y == 44 && x == 75)) oled_data <= 16'h2104;
            else if ((y == 36 && x == 67) || (y == 37 && x == 67) || (y == 29 && x == 68) || (y == 39 && x == 68) || (y == 29 && x == 69) || (y == 30 && x == 69) || (y == 39 && x == 69) || (y == 27 && x == 70) || (y == 28 && x == 70) || (y == 38 && x == 70) || (y == 39 && x == 70) || (y == 40 && x == 70) || (y == 41 && x == 70) || (y == 23 && x == 71) || (y == 27 && x == 71) || (y == 35 && x == 71) || (y == 36 && x == 71) || (y == 37 && x == 71) || (y == 38 && x == 71) || (y == 39 && x == 71) || (y == 40 && x == 71) || (y == 41 && x == 71) || (y == 25 && x == 72) || (y == 26 && x == 72) || (y == 37 && x == 72) || (y == 38 && x == 72) || (y == 39 && x == 72) || (y == 40 && x == 72) || (y == 41 && x == 72) || (y == 42 && x == 72) || (y == 43 && x == 72) || (y == 25 && x == 73) || (y == 26 && x == 73) || (y == 37 && x == 73) || (y == 38 && x == 73) || (y == 39 && x == 73) || (y == 40 && x == 73) || (y == 41 && x == 73) || (y == 42 && x == 73) || (y == 43 && x == 73) || (y == 23 && x == 74) || (y == 25 && x == 74) || (y == 26 && x == 74) || (y == 37 && x == 74) || (y == 38 && x == 74) || (y == 39 && x == 74) || (y == 40 && x == 74) || (y == 41 && x == 74) || (y == 42 && x == 74) || (y == 43 && x == 74) || (y == 23 && x == 75) || (y == 25 && x == 75) || (y == 26 && x == 75) || (y == 37 && x == 75) || (y == 38 && x == 75) || (y == 39 && x == 75) || (y == 40 && x == 75) || (y == 41 && x == 75) || (y == 42 && x == 75) || (y == 43 && x == 75) || (y == 24 && x == 76) || (y == 25 && x == 76) || (y == 26 && x == 76) || (y == 39 && x == 76) || (y == 40 && x == 76) || (y == 41 && x == 76) || (y == 42 && x == 76) || (y == 43 && x == 76) || (y == 24 && x == 77) || (y == 25 && x == 77) || (y == 26 && x == 77) || (y == 39 && x == 77) || (y == 40 && x == 77) || (y == 41 && x == 77) || (y == 23 && x == 78) || (y == 24 && x == 78) || (y == 25 && x == 78) || (y == 26 && x == 78) || (y == 27 && x == 78) || (y == 28 && x == 78) || (y == 35 && x == 78) || (y == 36 && x == 78) || (y == 37 && x == 78) || (y == 38 && x == 78) || (y == 39 && x == 78) || (y == 40 && x == 78) || (y == 41 && x == 78) || (y == 23 && x == 79) || (y == 25 && x == 79) || (y == 26 && x == 79) || (y == 27 && x == 79) || (y == 28 && x == 79) || (y == 35 && x == 79) || (y == 36 && x == 79) || (y == 37 && x == 79) || (y == 38 && x == 79) || (y == 39 && x == 79) || (y == 40 && x == 79) || (y == 41 && x == 79) || (y == 25 && x == 80) || (y == 26 && x == 80) || (y == 27 && x == 80) || (y == 28 && x == 80) || (y == 29 && x == 80) || (y == 30 && x == 80) || (y == 31 && x == 80) || (y == 32 && x == 80) || (y == 33 && x == 80) || (y == 34 && x == 80) || (y == 35 && x == 80) || (y == 36 && x == 80) || (y == 37 && x == 80) || (y == 38 && x == 80) || (y == 39 && x == 80) || (y == 40 && x == 80) || (y == 41 && x == 80) || (y == 27 && x == 81) || (y == 28 && x == 81) || (y == 29 && x == 81) || (y == 30 && x == 81) || (y == 31 && x == 81) || (y == 32 && x == 81) || (y == 33 && x == 81) || (y == 34 && x == 81) || (y == 35 && x == 81) || (y == 36 && x == 81) || (y == 37 && x == 81) || (y == 38 && x == 81) || (y == 39 && x == 81) || (y == 40 && x == 81) || (y == 41 && x == 81) || (y == 23 && x == 82) || (y == 27 && x == 82) || (y == 28 && x == 82) || (y == 29 && x == 82) || (y == 30 && x == 82) || (y == 31 && x == 82) || (y == 32 && x == 82) || (y == 33 && x == 82) || (y == 34 && x == 82) || (y == 35 && x == 82) || (y == 36 && x == 82) || (y == 37 && x == 82) || (y == 38 && x == 82) || (y == 39 && x == 82) || (y == 40 && x == 82) || (y == 41 && x == 82) || (y == 27 && x == 83) || (y == 28 && x == 83) || (y == 29 && x == 83) || (y == 30 && x == 83) || (y == 31 && x == 83) || (y == 32 && x == 83) || (y == 33 && x == 83) || (y == 34 && x == 83) || (y == 35 && x == 83) || (y == 36 && x == 83) || (y == 37 && x == 83) || (y == 38 && x == 83) || (y == 39 && x == 83) || (y == 27 && x == 84) || (y == 28 && x == 84) || (y == 29 && x == 84) || (y == 30 && x == 84) || (y == 31 && x == 84) || (y == 32 && x == 84) || (y == 33 && x == 84) || (y == 34 && x == 84) || (y == 35 && x == 84) || (y == 36 && x == 84) || (y == 37 && x == 84) || (y == 38 && x == 84) || (y == 39 && x == 84) || (y == 31 && x == 85) || (y == 32 && x == 85) || (y == 33 && x == 85) || (y == 34 && x == 85) || (y == 35 && x == 85) || (y == 31 && x == 86) || (y == 32 && x == 86) || (y == 33 && x == 86) || (y == 34 && x == 86) || (y == 35 && x == 86)) oled_data <= 16'h39a7;
            else if ((y == 46 && x == 75) || (y == 47 && x == 75) || (y == 48 && x == 75) || (y == 49 && x == 75) || (y == 44 && x == 77) || (y == 45 && x == 77) || (y == 43 && x == 85)) oled_data <= 16'h5201;
            else if ((y == 47 && x == 73) || (y == 44 && x == 88) || (y == 33 && x == 94) || (y == 34 && x == 94) || (y == 35 && x == 94)) oled_data <= 16'h2900;
            else if ((y == 31 && x == 66) || (y == 32 && x == 66) || (y == 38 && x == 66) || (y == 39 && x == 66) || (y == 31 && x == 67) || (y == 32 && x == 67) || (y == 39 && x == 67) || (y == 27 && x == 68) || (y == 28 && x == 68) || (y == 40 && x == 68) || (y == 41 && x == 68) || (y == 42 && x == 68) || (y == 43 && x == 68) || (y == 27 && x == 69) || (y == 28 && x == 69) || (y == 41 && x == 69) || (y == 42 && x == 69) || (y == 43 && x == 69) || (y == 25 && x == 70) || (y == 26 && x == 70) || (y == 42 && x == 70) || (y == 43 && x == 70) || (y == 25 && x == 71) || (y == 26 && x == 71) || (y == 42 && x == 71) || (y == 43 && x == 71) || (y == 44 && x == 72) || (y == 44 && x == 73) || (y == 45 && x == 73) || (y == 24 && x == 74) || (y == 44 && x == 74) || (y == 24 && x == 75) || (y == 24 && x == 80) || (y == 25 && x == 82) || (y == 26 && x == 82) || (y == 25 && x == 83) || (y == 26 && x == 83) || (y == 25 && x == 84) || (y == 26 && x == 84) || (y == 41 && x == 84) || (y == 40 && x == 85) || (y == 41 && x == 85) || (y == 27 && x == 86) || (y == 28 && x == 86) || (y == 29 && x == 86) || (y == 30 && x == 86) || (y == 37 && x == 86) || (y == 38 && x == 86) || (y == 39 && x == 86) || (y == 40 && x == 86) || (y == 41 && x == 86) || (y == 31 && x == 87) || (y == 32 && x == 87) || (y == 33 && x == 87) || (y == 34 && x == 87) || (y == 35 && x == 87) || (y == 36 && x == 87) || (y == 37 && x == 87) || (y == 31 && x == 88) || (y == 32 && x == 88) || (y == 33 && x == 88) || (y == 34 && x == 88) || (y == 35 && x == 88) || (y == 36 && x == 88) || (y == 37 && x == 88)) oled_data <= 16'h20e5;
            else if ((y == 46 && x == 86) || (y == 47 && x == 86) || (y == 33 && x == 91) || (y == 34 && x == 91) || (y == 35 && x == 91) || (y == 33 && x == 92) || (y == 34 && x == 92) || (y == 35 && x == 92)) oled_data <= 16'hdd87;
            else if ((y == 15 && x == 82)) oled_data <= 16'hfe03;
            else if ((y == 15 && x == 79) || (y == 16 && x == 81)) oled_data <= 16'hf520;
            else if ((y == 30 && x == 93) || (y == 30 && x == 94)) oled_data <= 16'hef39;
            else if ((y == 36 && x == 70) || (y == 37 && x == 70) || (y == 23 && x == 80) || (y == 25 && x == 81) || (y == 26 && x == 81) || (y == 40 && x == 83) || (y == 36 && x == 85) || (y == 36 && x == 86)) oled_data <= 16'h3146;
            else if ((y == 15 && x == 81)) oled_data <= 16'hfe64;
            else if ((y == 31 && x == 64) || (y == 32 && x == 64) || (y == 33 && x == 64) || (y == 34 && x == 64) || (y == 35 && x == 64) || (y == 36 && x == 64) || (y == 37 && x == 64) || (y == 38 && x == 64) || (y == 39 && x == 64) || (y == 21 && x == 74) || (y == 21 && x == 75)) oled_data <= 16'h7bef;
            else if ((y == 19 && x == 81)) oled_data <= 16'h834d;
            else if ((y == 37 && x == 69) || (y == 22 && x == 76) || (y == 37 && x == 76) || (y == 22 && x == 77) || (y == 36 && x == 77) || (y == 22 && x == 81) || (y == 21 && x == 82) || (y == 20 && x == 83)) oled_data <= 16'hce59;
            else if ((y == 15 && x == 77) || (y == 13 && x == 79)) oled_data <= 16'hfe53;
            else if ((y == 13 && x == 80) || (y == 13 && x == 81) || (y == 13 && x == 82)) oled_data <= 16'heb00;
            else if ((y == 34 && x == 71) || (y == 21 && x == 78) || (y == 34 && x == 78) || (y == 21 && x == 79) || (y == 29 && x == 79) || (y == 30 && x == 79) || (y == 31 && x == 79) || (y == 32 && x == 79) || (y == 33 && x == 79) || (y == 21 && x == 80) || (y == 22 && x == 83)) oled_data <= 16'h630d;
            else if ((y == 19 && x == 75)) oled_data <= 16'ha491;
            else if ((y == 48 && x == 79) || (y == 48 && x == 83)) oled_data <= 16'hd5a4;
            else if ((y == 36 && x == 93) || (y == 36 && x == 94)) oled_data <= 16'hb573;
            else if ((y == 44 && x == 79) || (y == 45 && x == 79) || (y == 49 && x == 79) || (y == 49 && x == 83)) oled_data <= 16'hc565;
            else if ((y == 48 && x == 69) || (y == 48 && x == 76) || (y == 49 && x == 77) || (y == 44 && x == 78) || (y == 45 && x == 78) || (y == 43 && x == 82) || (y == 43 && x == 83) || (y == 43 && x == 84) || (y == 49 && x == 85) || (y == 48 && x == 86) || (y == 30 && x == 92) || (y == 31 && x == 93) || (y == 31 && x == 94)) oled_data <= 16'hb4a6;
            else if ((y == 49 && x == 88)) oled_data <= 16'h4a04;
            else if ((y == 15 && x == 76) || (y == 14 && x == 77) || (y == 17 && x == 83) || (y == 14 && x == 85)) oled_data <= 16'hfef8;
            else if ((y == 12 && x == 79) || (y == 12 && x == 83) || (y == 13 && x == 83) || (y == 16 && x == 83)) oled_data <= 16'hfe75;
            else if ((y == 47 && x == 72)) oled_data <= 16'h20a0;
            else if ((y == 29 && x == 72) || (y == 30 && x == 72) || (y == 31 && x == 72) || (y == 32 && x == 72) || (y == 29 && x == 73) || (y == 30 && x == 73) || (y == 31 && x == 73) || (y == 32 && x == 73) || (y == 22 && x == 74) || (y == 29 && x == 74) || (y == 30 && x == 74) || (y == 31 && x == 74) || (y == 32 && x == 74) || (y == 22 && x == 75) || (y == 29 && x == 75) || (y == 30 && x == 75) || (y == 31 && x == 75) || (y == 32 && x == 75) || (y == 21 && x == 76) || (y == 21 && x == 81)) oled_data <= 16'h94f3;
            else if ((y == 44 && x == 85) || (y == 45 && x == 85)) oled_data <= 16'h5a61;
            else if ((y == 49 && x == 66)) oled_data <= 16'h6b0a;
            else if ((y == 47 && x == 67) || (y == 48 && x == 67) || (y == 50 && x == 69) || (y == 50 && x == 70) || (y == 50 && x == 71) || (y == 50 && x == 72) || (y == 50 && x == 73) || (y == 46 && x == 74) || (y == 47 && x == 74) || (y == 50 && x == 74) || (y == 50 && x == 75) || (y == 44 && x == 76) || (y == 50 && x == 76) || (y == 50 && x == 77) || (y == 42 && x == 78) || (y == 43 && x == 78) || (y == 50 && x == 78) || (y == 42 && x == 79) || (y == 50 && x == 79) || (y == 42 && x == 80) || (y == 50 && x == 80) || (y == 50 && x == 81) || (y == 50 && x == 82) || (y == 50 && x == 83) || (y == 50 && x == 84) || (y == 50 && x == 85) || (y == 42 && x == 86) || (y == 43 && x == 86) || (y == 44 && x == 86) || (y == 50 && x == 86) || (y == 45 && x == 87) || (y == 37 && x == 91) || (y == 37 && x == 92) || (y == 33 && x == 93) || (y == 34 && x == 93) || (y == 35 && x == 93)) oled_data <= 16'h39a2;
            else if ((y == 47 && x == 69) || (y == 47 && x == 76) || (y == 47 && x == 77) || (y == 47 && x == 78) || (y == 47 && x == 79) || (y == 44 && x == 80) || (y == 44 && x == 81) || (y == 44 && x == 83) || (y == 47 && x == 83) || (y == 47 && x == 84) || (y == 31 && x == 91) || (y == 32 && x == 91) || (y == 31 && x == 92)) oled_data <= 16'hfec6;
            else if ((y == 16 && x == 77) || (y == 17 && x == 77)) oled_data <= 16'hec03;
            else if ((y == 33 && x == 66) || (y == 34 && x == 66) || (y == 35 && x == 66) || (y == 36 && x == 66) || (y == 37 && x == 66) || (y == 33 && x == 67) || (y == 34 && x == 67) || (y == 35 && x == 67) || (y == 30 && x == 68) || (y == 28 && x == 71) || (y == 24 && x == 79) || (y == 23 && x == 81)) oled_data <= 16'h3166;
            else if ((y == 46 && x == 69) || (y == 46 && x == 70) || (y == 47 && x == 70) || (y == 48 && x == 70) || (y == 46 && x == 71) || (y == 47 && x == 71) || (y == 48 && x == 71) || (y == 48 && x == 72) || (y == 48 && x == 73) || (y == 46 && x == 76) || (y == 46 && x == 77) || (y == 16 && x == 78) || (y == 46 && x == 78) || (y == 16 && x == 79) || (y == 46 && x == 79) || (y == 14 && x == 80) || (y == 15 && x == 80) || (y == 16 && x == 80) || (y == 45 && x == 80) || (y == 46 && x == 80) || (y == 47 && x == 80) || (y == 48 && x == 80) || (y == 14 && x == 81) || (y == 45 && x == 81) || (y == 46 && x == 81) || (y == 47 && x == 81) || (y == 48 && x == 81) || (y == 14 && x == 82) || (y == 44 && x == 82) || (y == 45 && x == 82) || (y == 46 && x == 82) || (y == 47 && x == 82) || (y == 48 && x == 82) || (y == 45 && x == 83) || (y == 46 && x == 83) || (y == 44 && x == 84) || (y == 45 && x == 84) || (y == 46 && x == 84)) oled_data <= 16'hff05;
            else if ((y == 16 && x == 76) || (y == 17 && x == 76) || (y == 18 && x == 76) || (y == 18 && x == 77) || (y == 18 && x == 78) || (y == 18 && x == 79) || (y == 18 && x == 80)) oled_data <= 16'hf324;
            else if ((y == 38 && x == 67) || (y == 40 && x == 69) || (y == 35 && x == 70) || (y == 41 && x == 83) || (y == 40 && x == 84) || (y == 27 && x == 85) || (y == 28 && x == 85) || (y == 29 && x == 85) || (y == 30 && x == 85) || (y == 37 && x == 85) || (y == 38 && x == 85) || (y == 39 && x == 85)) oled_data <= 16'h2905;
            else if ((y == 19 && x == 74) || (y == 21 && x == 77) || (y == 19 && x == 82)) oled_data <= 16'h8c92;
            else if ((y == 19 && x == 76) || (y == 19 && x == 77) || (y == 19 && x == 78) || (y == 19 && x == 79) || (y == 19 && x == 80)) oled_data <= 16'h81e4;
            else if ((y == 37 && x == 68) || (y == 37 && x == 77)) oled_data <= 16'hb5b6;
            else if ((y == 44 && x == 66) || (y == 50 && x == 67) || (y == 24 && x == 69) || (y == 22 && x == 71) || (y == 20 && x == 73) || (y == 25 && x == 87) || (y == 26 && x == 88) || (y == 42 && x == 88) || (y == 43 && x == 88) || (y == 28 && x == 90) || (y == 37 && x == 93)) oled_data <= 16'hffdf;
            else if ((y == 14 && x == 79) || (y == 14 && x == 83)) oled_data <= 16'hf480;
            else if ((y == 14 && x == 78) || (y == 12 && x == 80) || (y == 12 && x == 81) || (y == 12 && x == 82) || (y == 16 && x == 82) || (y == 14 && x == 84)) oled_data <= 16'hf320;
            else if ((y == 48 && x == 74) || (y == 49 && x == 74) || (y == 45 && x == 76) || (y == 43 && x == 79) || (y == 43 && x == 80) || (y == 45 && x == 86) || (y == 46 && x == 87) || (y == 47 && x == 87) || (y == 48 && x == 87)) oled_data <= 16'h3940;
            else if ((y == 46 && x == 68) || (y == 32 && x == 92)) oled_data <= 16'hee88;
            else if ((y == 47 && x == 68) || (y == 49 && x == 70) || (y == 49 && x == 71) || (y == 49 && x == 72) || (y == 49 && x == 73) || (y == 49 && x == 80) || (y == 49 && x == 81) || (y == 49 && x == 82)) oled_data <= 16'hde26;
            else if ((y == 31 && x == 70) || (y == 32 && x == 70) || (y == 33 && x == 70) || (y == 27 && x == 77) || (y == 28 && x == 77) || (y == 21 && x == 83)) oled_data <= 16'h6b6e;
            else if ((y == 17 && x == 78) || (y == 17 && x == 79) || (y == 17 && x == 80)) oled_data <= 16'hfe07;
            else if ((y == 16 && x == 75) || (y == 17 && x == 75) || (y == 18 && x == 75) || (y == 15 && x == 85)) oled_data <= 16'hff5b;
            else if ((y == 46 && x == 66) || (y == 47 && x == 66) || (y == 48 && x == 66) || (y == 49 && x == 67) || (y == 50 && x == 68)) oled_data <= 16'h5246;
            else if ((y == 18 && x == 81)) oled_data <= 16'hf5d4;
            else if ((y == 43 && x == 81) || (y == 36 && x == 91) || (y == 36 && x == 92)) oled_data <= 16'h8363;
            else if ((y == 15 && x == 84)) oled_data <= 16'he428;
            else if ((y == 40 && x == 65) || (y == 36 && x == 68) || (y == 19 && x == 83) || (y == 21 && x == 85) || (y == 22 && x == 85) || (y == 23 && x == 85) || (y == 24 && x == 85) || (y == 38 && x == 89) || (y == 38 && x == 90)) oled_data <= 16'hd69a;
            else if ((y == 15 && x == 78)) oled_data <= 16'hf420;
            else if ((y == 42 && x == 81)) oled_data <= 16'h7305;
            else oled_data <= 16'hffff;
        end
        else if (count <= 150_000_000) begin
            if ((y == 28 && x == 66) || (y == 44 && x == 66) || (y == 24 && x == 83)) oled_data <= 16'h1062;
            else if ((y == 39 && x == 91) || (y == 39 && x == 92)) oled_data <= 16'hdeda;
            else if ((y == 22 && x == 72) || (y == 22 && x == 73) || (y == 22 && x == 84)) oled_data <= 16'h4a28;
            else if ((y == 18 && x == 82)) oled_data <= 16'hb34b;
            else if ((y == 47 && x == 67) || (y == 45 && x == 87) || (y == 46 && x == 88) || (y == 47 && x == 88) || (y == 48 && x == 88) || (y == 49 && x == 88)) oled_data <= 16'h3140;
            else if ((y == 30 && x == 91) || (y == 30 && x == 92)) oled_data <= 16'hb4a8;
            else if ((y == 23 && x == 83)) oled_data <= 16'h528a;
            else if ((y == 18 && x == 81)) oled_data <= 16'hf50c;
            else if ((y == 19 && x == 81)) oled_data <= 16'hcc70;
            else if ((y == 33 && x == 65) || (y == 34 && x == 65) || (y == 35 && x == 65) || (y == 36 && x == 65) || (y == 37 && x == 65) || (y == 38 && x == 65) || (y == 39 && x == 65) || (y == 29 && x == 67) || (y == 30 && x == 67) || (y == 42 && x == 67) || (y == 43 && x == 67) || (y == 26 && x == 68) || (y == 36 && x == 69) || (y == 36 && x == 70) || (y == 25 && x == 71) || (y == 21 && x == 75) || (y == 21 && x == 76) || (y == 36 && x == 76) || (y == 21 && x == 77) || (y == 36 && x == 77) || (y == 21 && x == 78) || (y == 36 && x == 78) || (y == 21 && x == 79) || (y == 21 && x == 80) || (y == 21 && x == 81) || (y == 21 && x == 82) || (y == 25 && x == 82) || (y == 25 && x == 83) || (y == 30 && x == 88) || (y == 31 && x == 89) || (y == 38 && x == 90)) oled_data <= 16'h841;
            else if ((y == 32 && x == 67) || (y == 40 && x == 67) || (y == 29 && x == 69) || (y == 41 && x == 69) || (y == 42 && x == 69) || (y == 43 && x == 69) || (y == 43 && x == 70) || (y == 27 && x == 71) || (y == 43 && x == 71) || (y == 45 && x == 72) || (y == 45 && x == 73) || (y == 45 && x == 74) || (y == 25 && x == 75) || (y == 25 && x == 80) || (y == 27 && x == 82) || (y == 27 && x == 83) || (y == 42 && x == 83) || (y == 27 && x == 84) || (y == 41 && x == 84) || (y == 42 && x == 84) || (y == 28 && x == 85) || (y == 29 && x == 85) || (y == 30 && x == 85) || (y == 38 && x == 85) || (y == 39 && x == 85) || (y == 40 && x == 85) || (y == 41 && x == 85) || (y == 42 && x == 85) || (y == 29 && x == 86) || (y == 30 && x == 86) || (y == 31 && x == 86) || (y == 38 && x == 86) || (y == 39 && x == 86) || (y == 40 && x == 86) || (y == 41 && x == 86) || (y == 42 && x == 86) || (y == 32 && x == 87) || (y == 33 && x == 87) || (y == 34 && x == 87) || (y == 35 && x == 87) || (y == 36 && x == 87) || (y == 37 && x == 87) || (y == 38 && x == 87) || (y == 33 && x == 88) || (y == 34 && x == 88) || (y == 35 && x == 88) || (y == 36 && x == 88) || (y == 38 && x == 88)) oled_data <= 16'hb122;
            else if ((y == 49 && x == 78) || (y == 49 && x == 79) || (y == 49 && x == 83) || (y == 49 && x == 84) || (y == 47 && x == 85) || (y == 48 && x == 85)) oled_data <= 16'hdd85;
            else if ((y == 17 && x == 75) || (y == 18 && x == 75) || (y == 19 && x == 75) || (y == 16 && x == 76) || (y == 15 && x == 77) || (y == 18 && x == 83) || (y == 15 && x == 85) || (y == 16 && x == 85)) oled_data <= 16'hff3b;
            else if ((y == 18 && x == 79)) oled_data <= 16'hebe6;
            else if ((y == 32 && x == 65) || (y == 40 && x == 65) || (y == 28 && x == 67) || (y == 44 && x == 67) || (y == 26 && x == 69) || (y == 27 && x == 69) || (y == 46 && x == 69) || (y == 25 && x == 70) || (y == 46 && x == 70) || (y == 36 && x == 71) || (y == 46 && x == 71) || (y == 23 && x == 72) || (y == 25 && x == 72) || (y == 47 && x == 72) || (y == 23 && x == 73) || (y == 25 && x == 73) || (y == 21 && x == 74) || (y == 25 && x == 84) || (y == 26 && x == 86) || (y == 27 && x == 86) || (y == 28 && x == 87) || (y == 28 && x == 88) || (y == 29 && x == 88) || (y == 40 && x == 88) || (y == 41 && x == 88) || (y == 42 && x == 88) || (y == 30 && x == 89) || (y == 30 && x == 90) || (y == 31 && x == 90) || (y == 32 && x == 90) || (y == 33 && x == 90) || (y == 34 && x == 90) || (y == 35 && x == 90) || (y == 36 && x == 90) || (y == 37 && x == 90) || (y == 30 && x == 95) || (y == 34 && x == 95) || (y == 36 && x == 95)) oled_data <= 16'h0;
            else if ((y == 49 && x == 77) || (y == 50 && x == 78) || (y == 50 && x == 84) || (y == 49 && x == 85) || (y == 31 && x == 91)) oled_data <= 16'hc4e6;
            else if ((y == 52 && x == 68) || (y == 52 && x == 69) || (y == 52 && x == 70) || (y == 52 && x == 71) || (y == 52 && x == 72) || (y == 52 && x == 73) || (y == 52 && x == 74) || (y == 52 && x == 75) || (y == 52 && x == 76) || (y == 52 && x == 77) || (y == 52 && x == 78) || (y == 52 && x == 79) || (y == 52 && x == 80) || (y == 52 && x == 81) || (y == 52 && x == 82) || (y == 52 && x == 83) || (y == 52 && x == 84) || (y == 52 && x == 85) || (y == 52 && x == 86)) oled_data <= 16'h9490;
            else if ((y == 36 && x == 72) || (y == 35 && x == 75) || (y == 37 && x == 75)) oled_data <= 16'he2c9;
            else if ((y == 20 && x == 77) || (y == 20 && x == 78) || (y == 20 && x == 79) || (y == 20 && x == 80)) oled_data <= 16'h7123;
            else if ((y == 17 && x == 81)) oled_data <= 16'hec85;
            else if ((y == 45 && x == 71) || (y == 24 && x == 72) || (y == 24 && x == 73) || (y == 47 && x == 73) || (y == 23 && x == 84) || (y == 24 && x == 84) || (y == 42 && x == 87)) oled_data <= 16'h800;
            else if ((y == 50 && x == 64) || (y == 46 && x == 66) || (y == 16 && x == 75) || (y == 14 && x == 78) || (y == 14 && x == 84) || (y == 51 && x == 87) || (y == 52 && x == 87) || (y == 45 && x == 89) || (y == 46 && x == 89) || (y == 47 && x == 89) || (y == 48 && x == 89) || (y == 49 && x == 89) || (y == 50 && x == 89)) oled_data <= 16'hffde;
            else if ((y == 31 && x == 68) || (y == 28 && x == 69) || (y == 44 && x == 69) || (y == 27 && x == 70) || (y == 44 && x == 70) || (y == 26 && x == 71) || (y == 44 && x == 71) || (y == 25 && x == 74) || (y == 46 && x == 74) || (y == 43 && x == 77) || (y == 26 && x == 82) || (y == 26 && x == 83) || (y == 26 && x == 84) || (y == 28 && x == 86) || (y == 32 && x == 88) || (y == 37 && x == 88)) oled_data <= 16'ha963;
            else if ((y == 36 && x == 79) || (y == 39 && x == 87)) oled_data <= 16'h48a2;
            else if ((y == 50 && x == 87)) oled_data <= 16'h5a64;
            else if ((y == 49 && x == 68) || (y == 50 && x == 68) || (y == 50 && x == 69) || (y == 50 && x == 76) || (y == 50 && x == 86) || (y == 33 && x == 93) || (y == 33 && x == 94)) oled_data <= 16'ha447;
            else if ((y == 39 && x == 88)) oled_data <= 16'h3881;
            else if ((y == 33 && x == 67) || (y == 39 && x == 67) || (y == 25 && x == 79) || (y == 26 && x == 81) || (y == 27 && x == 81) || (y == 41 && x == 83) || (y == 31 && x == 85) || (y == 37 && x == 85) || (y == 37 && x == 86)) oled_data <= 16'hc983;
            else if ((y == 17 && x == 79)) oled_data <= 16'hf466;
            else if ((y == 31 && x == 64) || (y == 41 && x == 64) || (y == 31 && x == 65)) oled_data <= 16'hef7d;
            else if ((y == 46 && x == 68)) oled_data <= 16'h20e3;
            else if ((y == 23 && x == 78) || (y == 23 && x == 79) || (y == 23 && x == 80)) oled_data <= 16'h73af;
            else if ((y == 13 && x == 79) || (y == 14 && x == 79) || (y == 13 && x == 83) || (y == 14 && x == 83) || (y == 17 && x == 83)) oled_data <= 16'he5d5;
            else if ((y == 16 && x == 84)) oled_data <= 16'hb2e9;
            else if ((y == 29 && x == 66) || (y == 30 && x == 66) || (y == 42 && x == 66) || (y == 43 && x == 66) || (y == 27 && x == 68) || (y == 45 && x == 68) || (y == 24 && x == 70)) oled_data <= 16'h2104;
            else if ((y == 24 && x == 71) || (y == 24 && x == 82)) oled_data <= 16'h39a7;
            else if ((y == 28 && x == 68) || (y == 29 && x == 68) || (y == 37 && x == 68) || (y == 41 && x == 68) || (y == 42 && x == 68) || (y == 43 && x == 68) || (y == 44 && x == 68) || (y == 26 && x == 70) || (y == 46 && x == 72) || (y == 46 && x == 73) || (y == 45 && x == 75) || (y == 46 && x == 75) || (y == 37 && x == 79)) oled_data <= 16'h9943;
            else if ((y == 47 && x == 75) || (y == 48 && x == 75) || (y == 49 && x == 75) || (y == 50 && x == 75) || (y == 45 && x == 77) || (y == 46 && x == 77) || (y == 44 && x == 85)) oled_data <= 16'h5201;
            else if ((y == 48 && x == 73) || (y == 45 && x == 88) || (y == 34 && x == 94) || (y == 35 && x == 94) || (y == 36 && x == 94)) oled_data <= 16'h2900;
            else if ((y == 18 && x == 80) || (y == 15 && x == 81) || (y == 16 && x == 81)) oled_data <= 16'hf546;
            else if ((y == 30 && x == 72) || (y == 31 && x == 72) || (y == 32 && x == 72) || (y == 30 && x == 73) || (y == 31 && x == 73) || (y == 32 && x == 73) || (y == 30 && x == 74) || (y == 31 && x == 74) || (y == 32 && x == 74)) oled_data <= 16'he3cf;
            else if ((y == 35 && x == 69) || (y == 35 && x == 70) || (y == 35 && x == 71) || (y == 24 && x == 74) || (y == 35 && x == 76) || (y == 35 && x == 77) || (y == 35 && x == 78)) oled_data <= 16'ha206;
            else if ((y == 47 && x == 86) || (y == 48 && x == 86) || (y == 34 && x == 91) || (y == 35 && x == 91) || (y == 36 && x == 91) || (y == 34 && x == 92) || (y == 35 && x == 92) || (y == 36 && x == 92)) oled_data <= 16'hdd87;
            else if ((y == 45 && x == 76) || (y == 43 && x == 78) || (y == 43 && x == 79) || (y == 43 && x == 80) || (y == 43 && x == 85) || (y == 43 && x == 86)) oled_data <= 16'h4161;
            else if ((y == 38 && x == 67) || (y == 38 && x == 69) || (y == 40 && x == 69) || (y == 38 && x == 70) || (y == 26 && x == 76) || (y == 27 && x == 76) || (y == 38 && x == 76) || (y == 38 && x == 78) || (y == 39 && x == 79) || (y == 36 && x == 80) || (y == 40 && x == 83) || (y == 28 && x == 84) || (y == 29 && x == 84) || (y == 30 && x == 84) || (y == 37 && x == 84) || (y == 39 && x == 84)) oled_data <= 16'hd9a4;
            else if ((y == 26 && x == 72) || (y == 37 && x == 72) || (y == 26 && x == 73) || (y == 37 && x == 73) || (y == 37 && x == 74) || (y == 30 && x == 79) || (y == 34 && x == 79)) oled_data <= 16'he226;
            else if ((y == 31 && x == 93) || (y == 31 && x == 94)) oled_data <= 16'hef39;
            else if ((y == 32 && x == 64) || (y == 33 && x == 64) || (y == 34 && x == 64) || (y == 35 && x == 64) || (y == 36 && x == 64) || (y == 37 && x == 64) || (y == 38 && x == 64) || (y == 39 && x == 64) || (y == 40 && x == 64) || (y == 22 && x == 74) || (y == 22 && x == 75)) oled_data <= 16'h7bef;
            else if ((y == 36 && x == 75) || (y == 24 && x == 76)) oled_data <= 16'hcac9;
            else if ((y == 20 && x == 81)) oled_data <= 16'h834d;
            else if ((y == 23 && x == 76) || (y == 23 && x == 81) || (y == 22 && x == 82) || (y == 21 && x == 83)) oled_data <= 16'hce59;
            else if ((y == 31 && x == 67) || (y == 41 && x == 67) || (y == 36 && x == 68) || (y == 27 && x == 85) || (y == 31 && x == 87) || (y == 31 && x == 88)) oled_data <= 16'h3041;
            else if ((y == 34 && x == 66) || (y == 35 && x == 66) || (y == 36 && x == 66) || (y == 37 && x == 66) || (y == 38 && x == 66) || (y == 35 && x == 68) || (y == 24 && x == 75) || (y == 24 && x == 80)) oled_data <= 16'ha9c5;
            else if ((y == 16 && x == 83)) oled_data <= 16'hc3a7;
            else if ((y == 43 && x == 82) || (y == 43 && x == 83) || (y == 43 && x == 84)) oled_data <= 16'hc487;
            else if ((y == 20 && x == 75)) oled_data <= 16'ha491;
            else if ((y == 22 && x == 78) || (y == 22 && x == 79) || (y == 22 && x == 80) || (y == 22 && x == 83)) oled_data <= 16'h630d;
            else if ((y == 37 && x == 93) || (y == 37 && x == 94)) oled_data <= 16'hb573;
            else if ((y == 45 && x == 79) || (y == 46 && x == 79) || (y == 50 && x == 79) || (y == 50 && x == 83)) oled_data <= 16'hc565;
            else if ((y == 30 && x == 68) || (y == 24 && x == 77) || (y == 24 && x == 78) || (y == 24 && x == 79) || (y == 35 && x == 79)) oled_data <= 16'hc227;
            else if ((y == 49 && x == 69) || (y == 49 && x == 76) || (y == 50 && x == 77) || (y == 45 && x == 78) || (y == 46 && x == 78) || (y == 44 && x == 82) || (y == 44 && x == 83) || (y == 44 && x == 84) || (y == 50 && x == 85) || (y == 49 && x == 86) || (y == 31 && x == 92) || (y == 32 && x == 93) || (y == 32 && x == 94)) oled_data <= 16'hb4a6;
            else if ((y == 47 && x == 66) || (y == 50 && x == 88)) oled_data <= 16'h4a04;
            else if ((y == 34 && x == 67) || (y == 35 && x == 67) || (y == 36 && x == 67) || (y == 37 && x == 67) || (y == 38 && x == 68) || (y == 39 && x == 68) || (y == 40 && x == 68) || (y == 30 && x == 69) || (y == 31 && x == 69) || (y == 39 && x == 69) || (y == 28 && x == 70) || (y == 29 && x == 70) || (y == 39 && x == 70) || (y == 40 && x == 70) || (y == 41 && x == 70) || (y == 42 && x == 70) || (y == 28 && x == 71) || (y == 29 && x == 71) || (y == 38 && x == 71) || (y == 39 && x == 71) || (y == 40 && x == 71) || (y == 41 && x == 71) || (y == 42 && x == 71) || (y == 27 && x == 72) || (y == 38 && x == 72) || (y == 39 && x == 72) || (y == 40 && x == 72) || (y == 41 && x == 72) || (y == 42 && x == 72) || (y == 43 && x == 72) || (y == 44 && x == 72) || (y == 27 && x == 73) || (y == 38 && x == 73) || (y == 39 && x == 73) || (y == 40 && x == 73) || (y == 41 && x == 73) || (y == 42 && x == 73) || (y == 43 && x == 73) || (y == 44 && x == 73) || (y == 26 && x == 74) || (y == 27 && x == 74) || (y == 38 && x == 74) || (y == 39 && x == 74) || (y == 40 && x == 74) || (y == 41 && x == 74) || (y == 42 && x == 74) || (y == 43 && x == 74) || (y == 44 && x == 74) || (y == 26 && x == 75) || (y == 27 && x == 75) || (y == 38 && x == 75) || (y == 39 && x == 75) || (y == 40 && x == 75) || (y == 41 && x == 75) || (y == 42 && x == 75) || (y == 43 && x == 75) || (y == 44 && x == 75) || (y == 25 && x == 76) || (y == 39 && x == 76) || (y == 40 && x == 76) || (y == 41 && x == 76) || (y == 42 && x == 76) || (y == 43 && x == 76) || (y == 44 && x == 76) || (y == 25 && x == 77) || (y == 26 && x == 77) || (y == 27 && x == 77) || (y == 38 && x == 77) || (y == 39 && x == 77) || (y == 40 && x == 77) || (y == 41 && x == 77) || (y == 42 && x == 77) || (y == 25 && x == 78) || (y == 26 && x == 78) || (y == 27 && x == 78) || (y == 28 && x == 78) || (y == 29 && x == 78) || (y == 39 && x == 78) || (y == 40 && x == 78) || (y == 41 && x == 78) || (y == 42 && x == 78) || (y == 26 && x == 79) || (y == 27 && x == 79) || (y == 28 && x == 79) || (y == 29 && x == 79) || (y == 38 && x == 79) || (y == 40 && x == 79) || (y == 41 && x == 79) || (y == 42 && x == 79) || (y == 26 && x == 80) || (y == 27 && x == 80) || (y == 28 && x == 80) || (y == 29 && x == 80) || (y == 30 && x == 80) || (y == 31 && x == 80) || (y == 32 && x == 80) || (y == 33 && x == 80) || (y == 34 && x == 80) || (y == 35 && x == 80) || (y == 37 && x == 80) || (y == 38 && x == 80) || (y == 39 && x == 80) || (y == 40 && x == 80) || (y == 41 && x == 80) || (y == 42 && x == 80) || (y == 28 && x == 81) || (y == 29 && x == 81) || (y == 30 && x == 81) || (y == 31 && x == 81) || (y == 32 && x == 81) || (y == 33 && x == 81) || (y == 34 && x == 81) || (y == 35 && x == 81) || (y == 36 && x == 81) || (y == 37 && x == 81) || (y == 38 && x == 81) || (y == 39 && x == 81) || (y == 40 && x == 81) || (y == 41 && x == 81) || (y == 42 && x == 81) || (y == 28 && x == 82) || (y == 29 && x == 82) || (y == 30 && x == 82) || (y == 31 && x == 82) || (y == 32 && x == 82) || (y == 33 && x == 82) || (y == 34 && x == 82) || (y == 35 && x == 82) || (y == 36 && x == 82) || (y == 37 && x == 82) || (y == 38 && x == 82) || (y == 39 && x == 82) || (y == 40 && x == 82) || (y == 41 && x == 82) || (y == 42 && x == 82) || (y == 28 && x == 83) || (y == 29 && x == 83) || (y == 30 && x == 83) || (y == 31 && x == 83) || (y == 32 && x == 83) || (y == 33 && x == 83) || (y == 34 && x == 83) || (y == 35 && x == 83) || (y == 36 && x == 83) || (y == 37 && x == 83) || (y == 38 && x == 83) || (y == 39 && x == 83) || (y == 31 && x == 84) || (y == 32 && x == 84) || (y == 33 && x == 84) || (y == 34 && x == 84) || (y == 35 && x == 84) || (y == 36 && x == 84) || (y == 38 && x == 84) || (y == 40 && x == 84) || (y == 32 && x == 85) || (y == 33 && x == 85) || (y == 34 && x == 85) || (y == 35 && x == 85) || (y == 36 && x == 85) || (y == 32 && x == 86) || (y == 33 && x == 86) || (y == 34 && x == 86) || (y == 35 && x == 86) || (y == 36 && x == 86)) oled_data <= 16'hd9c4;
            else if ((y == 48 && x == 72)) oled_data <= 16'h20a0;
            else if ((y == 23 && x == 74) || (y == 23 && x == 75) || (y == 22 && x == 76) || (y == 22 && x == 81)) oled_data <= 16'h94f3;
            else if ((y == 17 && x == 77) || (y == 18 && x == 77) || (y == 19 && x == 77) || (y == 16 && x == 78) || (y == 19 && x == 78) || (y == 15 && x == 79) || (y == 16 && x == 79)) oled_data <= 16'hca02;
            else if ((y == 33 && x == 72) || (y == 33 && x == 73) || (y == 33 && x == 74) || (y == 30 && x == 75) || (y == 31 && x == 75) || (y == 32 && x == 75) || (y == 33 && x == 75)) oled_data <= 16'heb6c;
            else if ((y == 45 && x == 85) || (y == 46 && x == 85)) oled_data <= 16'h5a61;
            else if ((y == 50 && x == 66)) oled_data <= 16'h6b0a;
            else if ((y == 48 && x == 67) || (y == 49 && x == 67) || (y == 51 && x == 69) || (y == 51 && x == 70) || (y == 51 && x == 71) || (y == 51 && x == 72) || (y == 51 && x == 73) || (y == 47 && x == 74) || (y == 48 && x == 74) || (y == 51 && x == 74) || (y == 51 && x == 75) || (y == 51 && x == 76) || (y == 51 && x == 77) || (y == 44 && x == 78) || (y == 51 && x == 78) || (y == 44 && x == 79) || (y == 51 && x == 79) || (y == 51 && x == 80) || (y == 51 && x == 81) || (y == 51 && x == 82) || (y == 51 && x == 83) || (y == 51 && x == 84) || (y == 51 && x == 85) || (y == 44 && x == 86) || (y == 45 && x == 86) || (y == 51 && x == 86) || (y == 46 && x == 87) || (y == 38 && x == 91) || (y == 38 && x == 92) || (y == 34 && x == 93) || (y == 35 && x == 93) || (y == 36 && x == 93)) oled_data <= 16'h39a2;
            else if ((y == 48 && x == 69) || (y == 48 && x == 76) || (y == 48 && x == 77) || (y == 48 && x == 78) || (y == 48 && x == 79) || (y == 45 && x == 80) || (y == 45 && x == 81) || (y == 48 && x == 83) || (y == 48 && x == 84) || (y == 32 && x == 91) || (y == 33 && x == 91) || (y == 32 && x == 92)) oled_data <= 16'hfec6;
            else if ((y == 16 && x == 80)) oled_data <= 16'hec03;
            else if ((y == 47 && x == 69) || (y == 47 && x == 70) || (y == 48 && x == 70) || (y == 49 && x == 70) || (y == 47 && x == 71) || (y == 48 && x == 71) || (y == 49 && x == 71) || (y == 49 && x == 72) || (y == 49 && x == 73) || (y == 47 && x == 76) || (y == 47 && x == 77) || (y == 47 && x == 78) || (y == 47 && x == 79) || (y == 17 && x == 80) || (y == 46 && x == 80) || (y == 47 && x == 80) || (y == 48 && x == 80) || (y == 49 && x == 80) || (y == 46 && x == 81) || (y == 47 && x == 81) || (y == 48 && x == 81) || (y == 49 && x == 81) || (y == 15 && x == 82) || (y == 45 && x == 82) || (y == 46 && x == 82) || (y == 47 && x == 82) || (y == 48 && x == 82) || (y == 49 && x == 82) || (y == 45 && x == 83) || (y == 46 && x == 83) || (y == 47 && x == 83) || (y == 45 && x == 84) || (y == 46 && x == 84) || (y == 47 && x == 84)) oled_data <= 16'hff05;
            else if ((y == 17 && x == 78) || (y == 18 && x == 78) || (y == 15 && x == 80)) oled_data <= 16'hf324;
            else if ((y == 20 && x == 74) || (y == 22 && x == 77) || (y == 20 && x == 82)) oled_data <= 16'h8c92;
            else if ((y == 23 && x == 77)) oled_data <= 16'hb5b6;
            else if ((y == 45 && x == 66) || (y == 51 && x == 67) || (y == 25 && x == 69) || (y == 23 && x == 70) || (y == 21 && x == 73) || (y == 12 && x == 80) || (y == 12 && x == 81) || (y == 12 && x == 82) || (y == 26 && x == 87) || (y == 27 && x == 88) || (y == 43 && x == 88) || (y == 44 && x == 88) || (y == 38 && x == 93)) oled_data <= 16'hffdf;
            else if ((y == 15 && x == 83)) oled_data <= 16'hc343;
            else if ((y == 44 && x == 77)) oled_data <= 16'hba86;
            else if ((y == 49 && x == 74) || (y == 50 && x == 74) || (y == 46 && x == 76) || (y == 44 && x == 80) || (y == 46 && x == 86) || (y == 47 && x == 87) || (y == 48 && x == 87) || (y == 49 && x == 87)) oled_data <= 16'h3940;
            else if ((y == 32 && x == 66) || (y == 33 && x == 66) || (y == 39 && x == 66) || (y == 40 && x == 66) || (y == 37 && x == 69) || (y == 37 && x == 70) || (y == 37 && x == 71) || (y == 37 && x == 76) || (y == 37 && x == 77) || (y == 37 && x == 78)) oled_data <= 16'h8944;
            else if ((y == 17 && x == 76) || (y == 18 && x == 76) || (y == 19 && x == 76) || (y == 15 && x == 78) || (y == 19 && x == 79) || (y == 13 && x == 80) || (y == 14 && x == 80) || (y == 19 && x == 80) || (y == 13 && x == 81) || (y == 14 && x == 81) || (y == 13 && x == 82) || (y == 14 && x == 82) || (y == 17 && x == 82) || (y == 15 && x == 84)) oled_data <= 16'hb940;
            else if ((y == 43 && x == 81)) oled_data <= 16'h8b25;
            else if ((y == 47 && x == 68) || (y == 33 && x == 92)) oled_data <= 16'hee88;
            else if ((y == 48 && x == 68) || (y == 50 && x == 70) || (y == 50 && x == 71) || (y == 50 && x == 72) || (y == 50 && x == 73) || (y == 50 && x == 80) || (y == 50 && x == 81) || (y == 50 && x == 82)) oled_data <= 16'hde26;
            else if ((y == 16 && x == 82)) oled_data <= 16'hfe07;
            else if ((y == 31 && x == 66) || (y == 41 && x == 66)) oled_data <= 16'h4124;
            else if ((y == 20 && x == 76) || (y == 25 && x == 81)) oled_data <= 16'h60a1;
            else if ((y == 48 && x == 66) || (y == 49 && x == 66) || (y == 50 && x == 67) || (y == 51 && x == 68)) oled_data <= 16'h5246;
            else if ((y == 16 && x == 77)) oled_data <= 16'hf5d4;
            else if ((y == 44 && x == 81) || (y == 37 && x == 91) || (y == 37 && x == 92)) oled_data <= 16'h8363;
            else if ((y == 32 && x == 68) || (y == 33 && x == 68) || (y == 34 && x == 68) || (y == 32 && x == 69) || (y == 33 && x == 69) || (y == 34 && x == 69) || (y == 30 && x == 70) || (y == 31 && x == 70) || (y == 32 && x == 70) || (y == 33 && x == 70) || (y == 34 && x == 70) || (y == 30 && x == 71) || (y == 31 && x == 71) || (y == 32 && x == 71) || (y == 33 && x == 71) || (y == 34 && x == 71) || (y == 28 && x == 72) || (y == 29 && x == 72) || (y == 34 && x == 72) || (y == 35 && x == 72) || (y == 28 && x == 73) || (y == 29 && x == 73) || (y == 34 && x == 73) || (y == 35 && x == 73) || (y == 36 && x == 73) || (y == 28 && x == 74) || (y == 29 && x == 74) || (y == 34 && x == 74) || (y == 35 && x == 74) || (y == 36 && x == 74) || (y == 28 && x == 75) || (y == 29 && x == 75) || (y == 34 && x == 75) || (y == 28 && x == 76) || (y == 29 && x == 76) || (y == 30 && x == 76) || (y == 31 && x == 76) || (y == 32 && x == 76) || (y == 33 && x == 76) || (y == 34 && x == 76) || (y == 28 && x == 77) || (y == 29 && x == 77) || (y == 30 && x == 77) || (y == 31 && x == 77) || (y == 32 && x == 77) || (y == 33 && x == 77) || (y == 34 && x == 77) || (y == 30 && x == 78) || (y == 31 && x == 78) || (y == 32 && x == 78) || (y == 33 && x == 78) || (y == 34 && x == 78) || (y == 31 && x == 79) || (y == 32 && x == 79) || (y == 33 && x == 79)) oled_data <= 16'heaa8;
            else if ((y == 24 && x == 81)) oled_data <= 16'h69c6;
            else if ((y == 41 && x == 65) || (y == 20 && x == 83) || (y == 22 && x == 85) || (y == 23 && x == 85) || (y == 24 && x == 85) || (y == 25 && x == 85) || (y == 39 && x == 89) || (y == 39 && x == 90)) oled_data <= 16'hd69a;
            else if ((y == 45 && x == 69) || (y == 45 && x == 70) || (y == 26 && x == 85) || (y == 29 && x == 87) || (y == 30 && x == 87) || (y == 40 && x == 87) || (y == 41 && x == 87) || (y == 32 && x == 89) || (y == 33 && x == 89) || (y == 34 && x == 89) || (y == 35 && x == 89) || (y == 36 && x == 89) || (y == 37 && x == 89) || (y == 38 && x == 89)) oled_data <= 16'h1800;
            else oled_data <= 16'hffff;
        end
        else if (count <= 200_000_000) begin
            if ((y == 48 && x == 75)) oled_data <= 16'h6980;
            else if ((y == 43 && x == 66)) oled_data <= 16'h1062;
            else if ((y == 44 && x == 66) || (y == 24 && x == 67) || (y == 44 && x == 67) || (y == 50 && x == 67)) oled_data <= 16'hffdf;
            else if ((y == 19 && x == 67) || (y == 19 && x == 68) || (y == 19 && x == 69) || (y == 19 && x == 70) || (y == 19 && x == 71) || (y == 19 && x == 72) || (y == 19 && x == 73) || (y == 19 && x == 74) || (y == 19 && x == 75) || (y == 19 && x == 76) || (y == 18 && x == 81) || (y == 19 && x == 82) || (y == 19 && x == 83) || (y == 19 && x == 84)) oled_data <= 16'he590;
            else if ((y == 16 && x == 79)) oled_data <= 16'hec8c;
            else if ((y == 32 && x == 94)) oled_data <= 16'hc3a7;
            else if ((y == 36 && x == 64) || (y == 37 && x == 66) || (y == 38 && x == 68) || (y == 38 && x == 69) || (y == 21 && x == 72) || (y == 21 && x == 73) || (y == 21 && x == 74) || (y == 23 && x == 77) || (y == 47 && x == 77) || (y == 41 && x == 79) || (y == 46 && x == 79) || (y == 47 && x == 79) || (y == 48 && x == 79) || (y == 21 && x == 81) || (y == 22 && x == 83) || (y == 38 && x == 83) || (y == 39 && x == 83) || (y == 42 && x == 83) || (y == 43 && x == 83) || (y == 44 && x == 83) || (y == 32 && x == 90) || (y == 32 && x == 91) || (y == 32 && x == 92) || (y == 36 && x == 92)) oled_data <= 16'hf480;
            else if ((y == 47 && x == 68)) oled_data <= 16'hc343;
            else if ((y == 48 && x == 68)) oled_data <= 16'h9c66;
            else if ((y == 48 && x == 74) || (y == 45 && x == 88) || (y == 46 && x == 88) || (y == 47 && x == 88) || (y == 48 && x == 88)) oled_data <= 16'h3140;
            else if ((y == 18 && x == 64) || (y == 19 && x == 64) || (y == 20 && x == 64) || (y == 25 && x == 64) || (y == 26 && x == 64) || (y == 39 && x == 64) || (y == 40 && x == 64) || (y == 41 && x == 64)) oled_data <= 16'he50d;
            else if ((y == 48 && x == 83)) oled_data <= 16'hd5a4;
            else if ((y == 29 && x == 79) || (y == 30 && x == 79)) oled_data <= 16'heef4;
            else if ((y == 49 && x == 83)) oled_data <= 16'hc565;
            else if ((y == 33 && x == 64) || (y == 18 && x == 65) || (y == 19 && x == 65) || (y == 20 && x == 65) || (y == 26 && x == 65) || (y == 33 && x == 65) || (y == 37 && x == 65) || (y == 38 && x == 65) || (y == 39 && x == 65) || (y == 40 && x == 65) || (y == 41 && x == 65) || (y == 20 && x == 66) || (y == 26 && x == 66) || (y == 39 && x == 66) || (y == 40 && x == 66) || (y == 41 && x == 66) || (y == 20 && x == 67) || (y == 21 && x == 67) || (y == 22 && x == 67) || (y == 26 && x == 67) || (y == 27 && x == 67) || (y == 28 && x == 67) || (y == 35 && x == 67) || (y == 39 && x == 67) || (y == 40 && x == 67) || (y == 41 && x == 67) || (y == 20 && x == 68) || (y == 21 && x == 68) || (y == 22 && x == 68) || (y == 25 && x == 68) || (y == 26 && x == 68) || (y == 27 && x == 68) || (y == 28 && x == 68) || (y == 20 && x == 69) || (y == 21 && x == 69) || (y == 22 && x == 69) || (y == 23 && x == 69) || (y == 24 && x == 69) || (y == 25 && x == 69) || (y == 26 && x == 69) || (y == 27 && x == 69) || (y == 28 && x == 69) || (y == 37 && x == 69) || (y == 46 && x == 69) || (y == 20 && x == 70) || (y == 21 && x == 70) || (y == 22 && x == 70) || (y == 25 && x == 70) || (y == 26 && x == 70) || (y == 43 && x == 70) || (y == 46 && x == 70) || (y == 47 && x == 70) || (y == 48 && x == 70) || (y == 20 && x == 71) || (y == 21 && x == 71) || (y == 22 && x == 71) || (y == 26 && x == 71) || (y == 42 && x == 71) || (y == 43 && x == 71) || (y == 46 && x == 71) || (y == 47 && x == 71) || (y == 48 && x == 71) || (y == 20 && x == 72) || (y == 44 && x == 72) || (y == 45 && x == 72) || (y == 46 && x == 72) || (y == 20 && x == 73) || (y == 45 && x == 73) || (y == 46 && x == 73) || (y == 20 && x == 74) || (y == 24 && x == 74) || (y == 20 && x == 75) || (y == 20 && x == 76) || (y == 21 && x == 76) || (y == 22 && x == 76) || (y == 25 && x == 76) || (y == 26 && x == 76) || (y == 48 && x == 76) || (y == 20 && x == 77) || (y == 21 && x == 77) || (y == 22 && x == 77) || (y == 48 && x == 77) || (y == 17 && x == 78) || (y == 18 && x == 78) || (y == 19 && x == 78) || (y == 20 && x == 78) || (y == 21 && x == 78) || (y == 22 && x == 78) || (y == 23 && x == 78) || (y == 24 && x == 78) || (y == 42 && x == 78) || (y == 43 && x == 78) || (y == 44 && x == 78) || (y == 45 && x == 78) || (y == 46 && x == 78) || (y == 47 && x == 78) || (y == 48 && x == 78) || (y == 18 && x == 79) || (y == 19 && x == 79) || (y == 20 && x == 79) || (y == 21 && x == 79) || (y == 22 && x == 79) || (y == 42 && x == 79) || (y == 43 && x == 79) || (y == 44 && x == 79) || (y == 45 && x == 79) || (y == 18 && x == 80) || (y == 19 && x == 80) || (y == 20 && x == 80) || (y == 21 && x == 80) || (y == 22 && x == 80) || (y == 41 && x == 80) || (y == 42 && x == 80) || (y == 43 && x == 80) || (y == 44 && x == 80) || (y == 20 && x == 81) || (y == 41 && x == 81) || (y == 42 && x == 81) || (y == 43 && x == 81) || (y == 44 && x == 81) || (y == 45 && x == 81) || (y == 20 && x == 82) || (y == 41 && x == 82) || (y == 42 && x == 82) || (y == 43 && x == 82) || (y == 44 && x == 82) || (y == 45 && x == 82) || (y == 46 && x == 82) || (y == 20 && x == 83) || (y == 40 && x == 83) || (y == 41 && x == 83) || (y == 20 && x == 84) || (y == 21 && x == 84) || (y == 22 && x == 84) || (y == 23 && x == 84) || (y == 24 && x == 84) || (y == 39 && x == 84) || (y == 40 && x == 84) || (y == 41 && x == 84) || (y == 24 && x == 85) || (y == 24 && x == 86) || (y == 27 && x == 86) || (y == 28 && x == 86) || (y == 43 && x == 86) || (y == 44 && x == 86) || (y == 24 && x == 87) || (y == 25 && x == 87) || (y == 26 && x == 87) || (y == 27 && x == 87) || (y == 28 && x == 87) || (y == 37 && x == 87) || (y == 25 && x == 88) || (y == 26 && x == 88) || (y == 27 && x == 88) || (y == 28 && x == 88) || (y == 29 && x == 88) || (y == 37 && x == 88) || (y == 41 && x == 88) || (y == 26 && x == 89) || (y == 27 && x == 89) || (y == 28 && x == 89) || (y == 29 && x == 89) || (y == 33 && x == 89) || (y == 37 && x == 89) || (y == 38 && x == 89) || (y == 39 && x == 89) || (y == 26 && x == 90) || (y == 33 && x == 90) || (y == 37 && x == 90) || (y == 38 && x == 90) || (y == 39 && x == 90) || (y == 26 && x == 91) || (y == 33 && x == 91) || (y == 37 && x == 91) || (y == 38 && x == 91) || (y == 39 && x == 91) || (y == 40 && x == 91) || (y == 41 && x == 91) || (y == 42 && x == 91) || (y == 42 && x == 92) || (y == 31 && x == 93)) oled_data <= 16'hf320;
            else if ((y == 48 && x == 69) || (y == 49 && x == 85) || (y == 48 && x == 86)) oled_data <= 16'hb4a6;
            else if ((y == 38 && x == 64) || (y == 19 && x == 66) || (y == 19 && x == 77)) oled_data <= 16'hf50c;
            else if ((y == 49 && x == 88)) oled_data <= 16'h4a04;
            else if ((y == 46 && x == 67) || (y == 49 && x == 74) || (y == 46 && x == 87) || (y == 47 && x == 87) || (y == 48 && x == 87)) oled_data <= 16'h3940;
            else if ((y == 32 && x == 65) || (y == 36 && x == 68) || (y == 39 && x == 68) || (y == 40 && x == 68) || (y == 41 && x == 68) || (y == 36 && x == 69) || (y == 23 && x == 70) || (y == 23 && x == 71) || (y == 22 && x == 75) || (y == 25 && x == 75) || (y == 26 && x == 75) || (y == 23 && x == 76) || (y == 47 && x == 76) || (y == 24 && x == 77) || (y == 42 && x == 77) || (y == 43 && x == 77) || (y == 46 && x == 77) || (y == 40 && x == 79) || (y == 23 && x == 80) || (y == 45 && x == 83) || (y == 38 && x == 85) || (y == 39 && x == 85) || (y == 40 && x == 85) || (y == 41 && x == 85) || (y == 38 && x == 87) || (y == 38 && x == 88) || (y == 32 && x == 89) || (y == 40 && x == 89) || (y == 40 && x == 90)) oled_data <= 16'hfce0;
            else if ((y == 23 && x == 68) || (y == 47 && x == 69) || (y == 27 && x == 90) || (y == 28 && x == 90) || (y == 29 && x == 90) || (y == 30 && x == 90) || (y == 25 && x == 92) || (y == 26 && x == 92) || (y == 33 && x == 92) || (y == 37 && x == 92) || (y == 38 && x == 92) || (y == 39 && x == 92) || (y == 40 && x == 92) || (y == 41 && x == 92) || (y == 42 && x == 93) || (y == 31 && x == 94) || (y == 43 && x == 94)) oled_data <= 16'heb62;
            else if ((y == 46 && x == 68) || (y == 49 && x == 70) || (y == 49 && x == 71) || (y == 49 && x == 76) || (y == 49 && x == 77) || (y == 49 && x == 78) || (y == 42 && x == 94)) oled_data <= 16'hcb21;
            else if ((y == 44 && x == 88)) oled_data <= 16'h2900;
            else if ((y == 44 && x == 87)) oled_data <= 16'h38c0;
            else if ((y == 35 && x == 66) || (y == 38 && x == 66) || (y == 38 && x == 67) || (y == 37 && x == 68) || (y == 42 && x == 70) || (y == 44 && x == 73) || (y == 23 && x == 74) || (y == 24 && x == 75) || (y == 25 && x == 77) || (y == 26 && x == 77) || (y == 40 && x == 80) || (y == 45 && x == 80) || (y == 40 && x == 81) || (y == 38 && x == 84) || (y == 27 && x == 85) || (y == 28 && x == 85) || (y == 42 && x == 85) || (y == 43 && x == 85) || (y == 44 && x == 85) || (y == 45 && x == 86) || (y == 40 && x == 87) || (y == 30 && x == 88) || (y == 40 && x == 88) || (y == 30 && x == 89)) oled_data <= 16'heb60;
            else if ((y == 42 && x == 68) || (y == 43 && x == 68) || (y == 44 && x == 68) || (y == 45 && x == 68) || (y == 47 && x == 74) || (y == 47 && x == 75) || (y == 30 && x == 80)) oled_data <= 16'hf546;
            else if ((y == 34 && x == 75) || (y == 37 && x == 75) || (y == 30 && x == 78) || (y == 30 && x == 91)) oled_data <= 16'hfffa;
            else if ((y == 17 && x == 64) || (y == 21 && x == 64) || (y == 18 && x == 66) || (y == 23 && x == 67) || (y == 16 && x == 77) || (y == 17 && x == 77) || (y == 18 && x == 77) || (y == 15 && x == 78) || (y == 20 && x == 85) || (y == 21 && x == 85) || (y == 22 && x == 85)) oled_data <= 16'hfef8;
            else if ((y == 48 && x == 84) || (y == 46 && x == 85) || (y == 47 && x == 85) || (y == 46 && x == 86)) oled_data <= 16'hdd85;
            else if ((y == 36 && x == 81)) oled_data <= 16'hee88;
            else if ((y == 29 && x == 64) || (y == 30 && x == 64) || (y == 31 && x == 64)) oled_data <= 16'hfeb0;
            else if ((y == 49 && x == 79)) oled_data <= 16'he446;
            else if ((y == 49 && x == 72) || (y == 49 && x == 73) || (y == 49 && x == 80) || (y == 49 && x == 81) || (y == 49 && x == 82)) oled_data <= 16'hde26;
            else if ((y == 47 && x == 86)) oled_data <= 16'hdd87;
            else if ((y == 21 && x == 65) || (y == 17 && x == 80)) oled_data <= 16'hfe75;
            else if ((y == 27 && x == 66) || (y == 28 && x == 66) || (y == 24 && x == 68) || (y == 17 && x == 79) || (y == 23 && x == 85) || (y == 23 && x == 86) || (y == 23 && x == 87) || (y == 23 && x == 88)) oled_data <= 16'hebe6;
            else if ((y == 32 && x == 64)) oled_data <= 16'hf5eb;
            else if ((y == 33 && x == 66) || (y == 38 && x == 77) || (y == 44 && x == 77) || (y == 45 && x == 77) || (y == 25 && x == 81) || (y == 26 && x == 81) || (y == 27 && x == 81) || (y == 28 && x == 81) || (y == 29 && x == 81) || (y == 37 && x == 81) || (y == 38 && x == 81) || (y == 39 && x == 81) || (y == 21 && x == 82) || (y == 36 && x == 82) || (y == 36 && x == 83) || (y == 46 && x == 83) || (y == 47 && x == 83) || (y == 36 && x == 84)) oled_data <= 16'hfe03;
            else if ((y == 17 && x == 66) || (y == 23 && x == 66) || (y == 17 && x == 81) || (y == 19 && x == 85) || (y == 30 && x == 93) || (y == 30 && x == 94)) oled_data <= 16'hff5b;
            else if ((y == 42 && x == 66)) oled_data <= 16'h20a0;
            else if ((y == 34 && x == 72) || (y == 32 && x == 74) || (y == 38 && x == 74) || (y == 29 && x == 77) || (y == 32 && x == 78)) oled_data <= 16'hf70d;
            else if ((y == 49 && x == 75) || (y == 45 && x == 87)) oled_data <= 16'h4161;
            else if ((y == 15 && x == 79)) oled_data <= 16'hff3b;
            else if ((y == 30 && x == 67) || (y == 34 && x == 67) || (y == 31 && x == 68) || (y == 32 && x == 68) || (y == 32 && x == 69) || (y == 40 && x == 70) || (y == 30 && x == 71) || (y == 40 && x == 71) || (y == 32 && x == 72) || (y == 32 && x == 73) || (y == 44 && x == 75) || (y == 38 && x == 76) || (y == 39 && x == 77) || (y == 40 && x == 78) || (y == 27 && x == 79) || (y == 28 && x == 79) || (y == 38 && x == 80) || (y == 23 && x == 82) || (y == 25 && x == 83) || (y == 26 && x == 83) || (y == 30 && x == 85) || (y == 35 && x == 85) || (y == 30 && x == 86)) oled_data <= 16'hed81;
            else if ((y == 42 && x == 67) || (y == 43 && x == 67)) oled_data <= 16'h0;
            else if ((y == 34 && x == 73) || (y == 30 && x == 77) || (y == 31 && x == 79)) oled_data <= 16'hff4f;
            else if ((y == 49 && x == 84) || (y == 48 && x == 85)) oled_data <= 16'hc4e6;
            else if ((y == 35 && x == 64) || (y == 29 && x == 65) || (y == 30 && x == 65) || (y == 31 && x == 65) || (y == 35 && x == 65) || (y == 29 && x == 66) || (y == 30 && x == 66) || (y == 34 && x == 66) || (y == 37 && x == 67) || (y == 30 && x == 68) || (y == 30 && x == 69) || (y == 31 && x == 69) || (y == 39 && x == 69) || (y == 40 && x == 69) || (y == 41 && x == 69) || (y == 42 && x == 69) || (y == 43 && x == 69) || (y == 44 && x == 69) || (y == 24 && x == 70) || (y == 29 && x == 70) || (y == 30 && x == 70) || (y == 35 && x == 70) || (y == 36 && x == 70) || (y == 41 && x == 70) || (y == 24 && x == 71) || (y == 27 && x == 71) || (y == 28 && x == 71) || (y == 29 && x == 71) || (y == 35 && x == 71) || (y == 36 && x == 71) || (y == 37 && x == 71) || (y == 41 && x == 71) || (y == 22 && x == 72) || (y == 23 && x == 72) || (y == 24 && x == 72) || (y == 31 && x == 72) || (y == 42 && x == 72) || (y == 22 && x == 73) || (y == 23 && x == 73) || (y == 31 && x == 73) || (y == 42 && x == 73) || (y == 43 && x == 73) || (y == 22 && x == 74) || (y == 25 && x == 74) || (y == 26 && x == 74) || (y == 44 && x == 74) || (y == 45 && x == 74) || (y == 45 && x == 75) || (y == 46 && x == 75) || (y == 24 && x == 76) || (y == 27 && x == 76) || (y == 28 && x == 76) || (y == 39 && x == 76) || (y == 42 && x == 76) || (y == 43 && x == 76) || (y == 46 && x == 76) || (y == 27 && x == 77) || (y == 28 && x == 77) || (y == 26 && x == 78) || (y == 27 && x == 78) || (y == 28 && x == 78) || (y == 41 && x == 78) || (y == 25 && x == 79) || (y == 26 && x == 79) || (y == 24 && x == 80) || (y == 25 && x == 80) || (y == 26 && x == 80) || (y == 29 && x == 80) || (y == 39 && x == 80) || (y == 22 && x == 81) || (y == 23 && x == 81) || (y == 24 && x == 81) || (y == 47 && x == 81) || (y == 24 && x == 82) || (y == 27 && x == 82) || (y == 28 && x == 82) || (y == 37 && x == 82) || (y == 27 && x == 83) || (y == 28 && x == 83) || (y == 37 && x == 83) || (y == 26 && x == 84) || (y == 27 && x == 84) || (y == 28 && x == 84) || (y == 37 && x == 84) || (y == 43 && x == 84) || (y == 44 && x == 84) || (y == 45 && x == 84) || (y == 26 && x == 85) || (y == 29 && x == 85) || (y == 36 && x == 85) || (y == 37 && x == 85) || (y == 26 && x == 86) || (y == 35 && x == 86) || (y == 36 && x == 86) || (y == 37 && x == 86) || (y == 38 && x == 86) || (y == 39 && x == 86) || (y == 40 && x == 86) || (y == 41 && x == 86) || (y == 33 && x == 87) || (y == 34 && x == 87) || (y == 35 && x == 87) || (y == 39 && x == 87) || (y == 34 && x == 88) || (y == 35 && x == 88) || (y == 39 && x == 88) || (y == 31 && x == 89) || (y == 35 && x == 89) || (y == 42 && x == 89) || (y == 43 && x == 89) || (y == 31 && x == 90) || (y == 35 && x == 90) || (y == 31 && x == 91) || (y == 35 && x == 91) || (y == 35 && x == 92)) oled_data <= 16'hf520;
            else if ((y == 49 && x == 66)) oled_data <= 16'h6b0a;
            else if ((y == 47 && x == 67) || (y == 48 && x == 67) || (y == 50 && x == 69) || (y == 50 && x == 70) || (y == 50 && x == 71) || (y == 50 && x == 72) || (y == 50 && x == 73) || (y == 50 && x == 74) || (y == 50 && x == 75) || (y == 50 && x == 76) || (y == 50 && x == 77) || (y == 50 && x == 78) || (y == 50 && x == 79) || (y == 50 && x == 80) || (y == 50 && x == 81) || (y == 50 && x == 82) || (y == 50 && x == 83) || (y == 50 && x == 84) || (y == 50 && x == 85) || (y == 50 && x == 86)) oled_data <= 16'h39a2;
            else if ((y == 51 && x == 68) || (y == 51 && x == 69) || (y == 51 && x == 70) || (y == 51 && x == 71) || (y == 51 && x == 72) || (y == 51 && x == 73) || (y == 51 && x == 74) || (y == 51 && x == 75) || (y == 51 && x == 76) || (y == 51 && x == 77) || (y == 51 && x == 78) || (y == 51 && x == 79) || (y == 51 && x == 80) || (y == 51 && x == 81) || (y == 51 && x == 82) || (y == 51 && x == 83) || (y == 51 && x == 84) || (y == 51 && x == 85) || (y == 51 && x == 86)) oled_data <= 16'h9490;
            else if ((y == 21 && x == 66) || (y == 30 && x == 87) || (y == 34 && x == 92)) oled_data <= 16'hec03;
            else if ((y == 46 && x == 66) || (y == 47 && x == 66) || (y == 48 && x == 66) || (y == 49 && x == 67) || (y == 50 && x == 68)) oled_data <= 16'h5246;
            else if ((y == 34 && x == 68) || (y == 30 && x == 72) || (y == 30 && x == 73) || (y == 33 && x == 73) || (y == 37 && x == 73) || (y == 35 && x == 74) || (y == 27 && x == 75) || (y == 28 && x == 75) || (y == 30 && x == 75) || (y == 39 && x == 75) || (y == 42 && x == 75) || (y == 43 && x == 75) || (y == 40 && x == 76) || (y == 47 && x == 84)) oled_data <= 16'hfec6;
            else if ((y == 22 && x == 66) || (y == 19 && x == 81) || (y == 32 && x == 93)) oled_data <= 16'he428;
            else if ((y == 29 && x == 67) || (y == 29 && x == 68) || (y == 29 && x == 69) || (y == 45 && x == 69) || (y == 27 && x == 70) || (y == 28 && x == 70) || (y == 37 && x == 70) || (y == 44 && x == 70) || (y == 45 && x == 70) || (y == 44 && x == 71) || (y == 45 && x == 71) || (y == 43 && x == 72) || (y == 24 && x == 73) || (y == 46 && x == 74) || (y == 25 && x == 78) || (y == 46 && x == 81) || (y == 25 && x == 84) || (y == 42 && x == 84) || (y == 25 && x == 85) || (y == 25 && x == 86) || (y == 29 && x == 86) || (y == 33 && x == 88) || (y == 41 && x == 89) || (y == 41 && x == 90) || (y == 42 && x == 90) || (y == 43 && x == 90) || (y == 31 && x == 92)) oled_data <= 16'hfd00;
            else if ((y == 31 && x == 75) || (y == 35 && x == 75) || (y == 38 && x == 75) || (y == 30 && x == 76)) oled_data <= 16'hff2a;
            else if ((y == 31 && x == 67) || (y == 32 && x == 67) || (y == 33 && x == 67) || (y == 33 && x == 68) || (y == 33 && x == 69) || (y == 34 && x == 69) || (y == 35 && x == 69) || (y == 31 && x == 70) || (y == 32 && x == 70) || (y == 33 && x == 70) || (y == 39 && x == 70) || (y == 31 && x == 71) || (y == 32 && x == 71) || (y == 33 && x == 71) || (y == 39 && x == 71) || (y == 25 && x == 72) || (y == 26 && x == 72) || (y == 27 && x == 72) || (y == 28 && x == 72) || (y == 29 && x == 72) || (y == 33 && x == 72) || (y == 37 && x == 72) || (y == 38 && x == 72) || (y == 39 && x == 72) || (y == 40 && x == 72) || (y == 41 && x == 72) || (y == 48 && x == 72) || (y == 25 && x == 73) || (y == 26 && x == 73) || (y == 27 && x == 73) || (y == 28 && x == 73) || (y == 29 && x == 73) || (y == 38 && x == 73) || (y == 39 && x == 73) || (y == 40 && x == 73) || (y == 41 && x == 73) || (y == 48 && x == 73) || (y == 27 && x == 74) || (y == 28 && x == 74) || (y == 29 && x == 74) || (y == 30 && x == 74) || (y == 31 && x == 74) || (y == 39 && x == 74) || (y == 40 && x == 74) || (y == 41 && x == 74) || (y == 42 && x == 74) || (y == 43 && x == 74) || (y == 29 && x == 75) || (y == 40 && x == 75) || (y == 41 && x == 75) || (y == 29 && x == 76) || (y == 37 && x == 76) || (y == 41 && x == 76) || (y == 44 && x == 76) || (y == 45 && x == 76) || (y == 37 && x == 77) || (y == 31 && x == 78) || (y == 37 && x == 78) || (y == 38 && x == 78) || (y == 39 && x == 78) || (y == 37 && x == 79) || (y == 27 && x == 80) || (y == 28 && x == 80) || (y == 37 && x == 80) || (y == 46 && x == 80) || (y == 47 && x == 80) || (y == 48 && x == 80) || (y == 48 && x == 81) || (y == 22 && x == 82) || (y == 25 && x == 82) || (y == 26 && x == 82) || (y == 29 && x == 82) || (y == 30 && x == 82) || (y == 31 && x == 82) || (y == 32 && x == 82) || (y == 33 && x == 82) || (y == 34 && x == 82) || (y == 35 && x == 82) || (y == 39 && x == 82) || (y == 48 && x == 82) || (y == 29 && x == 83) || (y == 30 && x == 83) || (y == 31 && x == 83) || (y == 32 && x == 83) || (y == 33 && x == 83) || (y == 34 && x == 83) || (y == 35 && x == 83) || (y == 29 && x == 84) || (y == 30 && x == 84) || (y == 31 && x == 84) || (y == 32 && x == 84) || (y == 33 && x == 84) || (y == 34 && x == 84) || (y == 35 && x == 84) || (y == 46 && x == 84) || (y == 31 && x == 85) || (y == 32 && x == 85) || (y == 33 && x == 85) || (y == 31 && x == 86) || (y == 32 && x == 86) || (y == 33 && x == 86) || (y == 31 && x == 87) || (y == 31 && x == 88)) oled_data <= 16'hff05;
            else if ((y == 42 && x == 88)) oled_data <= 16'hef39;
            else if ((y == 31 && x == 66) || (y == 32 && x == 66) || (y == 35 && x == 68) || (y == 34 && x == 70) || (y == 38 && x == 70) || (y == 34 && x == 71) || (y == 38 && x == 71) || (y == 40 && x == 77) || (y == 41 && x == 77) || (y == 38 && x == 79) || (y == 39 && x == 79) || (y == 30 && x == 81) || (y == 38 && x == 82) || (y == 34 && x == 85) || (y == 34 && x == 86) || (y == 32 && x == 87) || (y == 32 && x == 88)) oled_data <= 16'hfe64;
            else if ((y == 34 && x == 74) || (y == 31 && x == 77)) oled_data <= 16'hfff7;
            else if ((y == 27 && x == 64) || (y == 28 && x == 64) || (y == 45 && x == 66) || (y == 50 && x == 87) || (y == 51 && x == 87) || (y == 45 && x == 89) || (y == 46 && x == 89) || (y == 47 && x == 89) || (y == 48 && x == 89) || (y == 49 && x == 89) || (y == 28 && x == 91) || (y == 29 && x == 91) || (y == 27 && x == 92) || (y == 41 && x == 93) || (y == 41 && x == 94)) oled_data <= 16'hffde;
            else if ((y == 49 && x == 87)) oled_data <= 16'h5a64;
            else if ((y == 49 && x == 68) || (y == 49 && x == 69) || (y == 49 && x == 86)) oled_data <= 16'ha447;
            else if ((y == 16 && x == 78)) oled_data <= 16'hf324;
            else if ((y == 17 && x == 65)) oled_data <= 16'hfe53;
            else if ((y == 36 && x == 72) || (y == 36 && x == 73) || (y == 36 && x == 74) || (y == 32 && x == 75) || (y == 36 && x == 75) || (y == 36 && x == 76) || (y == 36 && x == 77) || (y == 36 && x == 78) || (y == 32 && x == 79) || (y == 36 && x == 79) || (y == 36 && x == 80) || (y == 31 && x == 81) || (y == 32 && x == 81) || (y == 33 && x == 81) || (y == 34 && x == 81) || (y == 35 && x == 81)) oled_data <= 16'hff72;
            else if ((y == 34 && x == 64) || (y == 34 && x == 65) || (y == 47 && x == 72) || (y == 47 && x == 73) || (y == 23 && x == 75) || (y == 23 && x == 79) || (y == 24 && x == 79) || (y == 40 && x == 82) || (y == 47 && x == 82) || (y == 21 && x == 83) || (y == 23 && x == 83) || (y == 24 && x == 83) || (y == 45 && x == 85) || (y == 34 && x == 89) || (y == 34 && x == 90) || (y == 34 && x == 91)) oled_data <= 16'hf3e0;
            else if ((y == 37 && x == 64) || (y == 36 && x == 65) || (y == 36 && x == 66) || (y == 36 && x == 67) || (y == 21 && x == 75) || (y == 36 && x == 87) || (y == 36 && x == 88) || (y == 36 && x == 89) || (y == 36 && x == 90) || (y == 36 && x == 91)) oled_data <= 16'hf420;
            else if ((y == 25 && x == 65) || (y == 25 && x == 66) || (y == 25 && x == 67) || (y == 25 && x == 71) || (y == 42 && x == 86) || (y == 29 && x == 87) || (y == 41 && x == 87) || (y == 24 && x == 88) || (y == 25 && x == 89) || (y == 25 && x == 90) || (y == 25 && x == 91) || (y == 43 && x == 91) || (y == 43 && x == 92) || (y == 43 && x == 93)) oled_data <= 16'heb00;
            else if ((y == 32 && x == 77) || (y == 42 && x == 87) || (y == 30 && x == 92)) oled_data <= 16'hffda;
            else if ((y == 42 && x == 64) || (y == 27 && x == 65) || (y == 28 && x == 65) || (y == 42 && x == 65) || (y == 15 && x == 77) || (y == 43 && x == 87) || (y == 23 && x == 89) || (y == 24 && x == 89) || (y == 44 && x == 89) || (y == 44 && x == 90) || (y == 27 && x == 91) || (y == 44 && x == 91) || (y == 44 && x == 92) || (y == 44 && x == 93) || (y == 44 && x == 94)) oled_data <= 16'hffbd;
            else oled_data <= 16'hffff;
        end
        else oled_data <= 16'hffff;
        count = (count == 200_000_000) ? 0 : count + 1;
    end
endmodule
